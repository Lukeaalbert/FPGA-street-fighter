module samurai_sprite
	(
		input wire clk,
		input wire [6:0] row,
		input wire [6:0] col,
		output reg [11:0] color_data
	);

	(* rom_style = "block" *)

	//signal declaration
	reg [6:0] row_reg;
	reg [6:0] col_reg;

	always @(posedge clk)
		begin
		row_reg <= row;
		col_reg <= col;
		end

	always @(*) begin

		if(({row_reg, col_reg}>=14'b00000000000000) && ({row_reg, col_reg}<14'b00000010110010)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=14'b00000010110010) && ({row_reg, col_reg}<14'b00000010110100)) color_data = 12'b000000001110;
		if(({row_reg, col_reg}>=14'b00000010110100) && ({row_reg, col_reg}<14'b00000010110111)) color_data = 12'b000000001101;
		if(({row_reg, col_reg}>=14'b00000010110111) && ({row_reg, col_reg}<14'b00000010111001)) color_data = 12'b000000001110;

		if(({row_reg, col_reg}>=14'b00000010111001) && ({row_reg, col_reg}<14'b00000100110001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==14'b00000100110001)) color_data = 12'b000000001110;
		if(({row_reg, col_reg}==14'b00000100110010)) color_data = 12'b000000001100;
		if(({row_reg, col_reg}==14'b00000100110011)) color_data = 12'b000000001011;
		if(({row_reg, col_reg}>=14'b00000100110100) && ({row_reg, col_reg}<14'b00000100110111)) color_data = 12'b000000001001;
		if(({row_reg, col_reg}==14'b00000100110111)) color_data = 12'b000000001010;
		if(({row_reg, col_reg}==14'b00000100111000)) color_data = 12'b000000001011;
		if(({row_reg, col_reg}==14'b00000100111001)) color_data = 12'b000000001101;
		if(({row_reg, col_reg}==14'b00000100111010)) color_data = 12'b000000001110;

		if(({row_reg, col_reg}>=14'b00000100111011) && ({row_reg, col_reg}<14'b00000110110000)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==14'b00000110110000)) color_data = 12'b000000001110;
		if(({row_reg, col_reg}==14'b00000110110001)) color_data = 12'b000000001100;
		if(({row_reg, col_reg}==14'b00000110110010)) color_data = 12'b000000001001;
		if(({row_reg, col_reg}==14'b00000110110011)) color_data = 12'b000000000111;
		if(({row_reg, col_reg}>=14'b00000110110100) && ({row_reg, col_reg}<14'b00000110110111)) color_data = 12'b000100000101;
		if(({row_reg, col_reg}==14'b00000110110111)) color_data = 12'b000000000110;
		if(({row_reg, col_reg}==14'b00000110111000)) color_data = 12'b000000001000;
		if(({row_reg, col_reg}==14'b00000110111001)) color_data = 12'b000000001010;
		if(({row_reg, col_reg}==14'b00000110111010)) color_data = 12'b000000001100;
		if(({row_reg, col_reg}==14'b00000110111011)) color_data = 12'b000000001101;
		if(({row_reg, col_reg}==14'b00000110111100)) color_data = 12'b000000001110;

		if(({row_reg, col_reg}>=14'b00000110111101) && ({row_reg, col_reg}<14'b00001000101111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==14'b00001000101111)) color_data = 12'b000000001110;
		if(({row_reg, col_reg}==14'b00001000110000)) color_data = 12'b000100001100;
		if(({row_reg, col_reg}==14'b00001000110001)) color_data = 12'b000100001010;
		if(({row_reg, col_reg}==14'b00001000110010)) color_data = 12'b000100000111;
		if(({row_reg, col_reg}==14'b00001000110011)) color_data = 12'b001100010101;
		if(({row_reg, col_reg}>=14'b00001000110100) && ({row_reg, col_reg}<14'b00001000110111)) color_data = 12'b010000100100;
		if(({row_reg, col_reg}==14'b00001000110111)) color_data = 12'b001100100101;
		if(({row_reg, col_reg}==14'b00001000111000)) color_data = 12'b000100000101;
		if(({row_reg, col_reg}==14'b00001000111001)) color_data = 12'b000100000111;
		if(({row_reg, col_reg}==14'b00001000111010)) color_data = 12'b000100001001;
		if(({row_reg, col_reg}==14'b00001000111011)) color_data = 12'b000000001010;
		if(({row_reg, col_reg}==14'b00001000111100)) color_data = 12'b000000001011;
		if(({row_reg, col_reg}==14'b00001000111101)) color_data = 12'b000000001101;

		if(({row_reg, col_reg}>=14'b00001000111110) && ({row_reg, col_reg}<14'b00001010101110)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=14'b00001010101110) && ({row_reg, col_reg}<14'b00001010110000)) color_data = 12'b000000001110;
		if(({row_reg, col_reg}==14'b00001010110000)) color_data = 12'b000000001001;
		if(({row_reg, col_reg}==14'b00001010110001)) color_data = 12'b000100001000;
		if(({row_reg, col_reg}==14'b00001010110010)) color_data = 12'b001000010101;
		if(({row_reg, col_reg}==14'b00001010110011)) color_data = 12'b010000100100;
		if(({row_reg, col_reg}==14'b00001010110100)) color_data = 12'b010100100011;
		if(({row_reg, col_reg}>=14'b00001010110101) && ({row_reg, col_reg}<14'b00001010110111)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}==14'b00001010110111)) color_data = 12'b010000100100;
		if(({row_reg, col_reg}==14'b00001010111000)) color_data = 12'b001100010100;
		if(({row_reg, col_reg}==14'b00001010111001)) color_data = 12'b001000010101;
		if(({row_reg, col_reg}==14'b00001010111010)) color_data = 12'b000100000110;
		if(({row_reg, col_reg}==14'b00001010111011)) color_data = 12'b000100000111;
		if(({row_reg, col_reg}==14'b00001010111100)) color_data = 12'b000000001000;
		if(({row_reg, col_reg}==14'b00001010111101)) color_data = 12'b000000001010;
		if(({row_reg, col_reg}==14'b00001010111110)) color_data = 12'b000000001100;
		if(({row_reg, col_reg}==14'b00001010111111)) color_data = 12'b000000001110;

		if(({row_reg, col_reg}>=14'b00001011000000) && ({row_reg, col_reg}<14'b00001100101110)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=14'b00001100101110) && ({row_reg, col_reg}<14'b00001100110000)) color_data = 12'b000000001110;
		if(({row_reg, col_reg}==14'b00001100110000)) color_data = 12'b000100000111;
		if(({row_reg, col_reg}==14'b00001100110001)) color_data = 12'b001100010111;
		if(({row_reg, col_reg}==14'b00001100110010)) color_data = 12'b010000100101;
		if(({row_reg, col_reg}==14'b00001100110011)) color_data = 12'b010000100011;
		if(({row_reg, col_reg}==14'b00001100110100)) color_data = 12'b010100100010;
		if(({row_reg, col_reg}>=14'b00001100110101) && ({row_reg, col_reg}<14'b00001100110111)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}==14'b00001100110111)) color_data = 12'b010000100011;
		if(({row_reg, col_reg}==14'b00001100111000)) color_data = 12'b010000100100;
		if(({row_reg, col_reg}>=14'b00001100111001) && ({row_reg, col_reg}<14'b00001100111011)) color_data = 12'b001100010100;
		if(({row_reg, col_reg}==14'b00001100111011)) color_data = 12'b001000010101;
		if(({row_reg, col_reg}==14'b00001100111100)) color_data = 12'b000100000101;
		if(({row_reg, col_reg}==14'b00001100111101)) color_data = 12'b000000000111;
		if(({row_reg, col_reg}==14'b00001100111110)) color_data = 12'b000000001001;
		if(({row_reg, col_reg}==14'b00001100111111)) color_data = 12'b000000001011;

		if(({row_reg, col_reg}>=14'b00001101000000) && ({row_reg, col_reg}<14'b00001110101110)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=14'b00001110101110) && ({row_reg, col_reg}<14'b00001110110000)) color_data = 12'b000000001110;
		if(({row_reg, col_reg}==14'b00001110110000)) color_data = 12'b000100000110;
		if(({row_reg, col_reg}==14'b00001110110001)) color_data = 12'b010000100110;
		if(({row_reg, col_reg}==14'b00001110110010)) color_data = 12'b010100100101;
		if(({row_reg, col_reg}>=14'b00001110110011) && ({row_reg, col_reg}<14'b00001110110101)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}==14'b00001110110101)) color_data = 12'b010100100010;
		if(({row_reg, col_reg}==14'b00001110110110)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}>=14'b00001110110111) && ({row_reg, col_reg}<14'b00001110111001)) color_data = 12'b010000100011;
		if(({row_reg, col_reg}==14'b00001110111001)) color_data = 12'b010000010011;
		if(({row_reg, col_reg}>=14'b00001110111010) && ({row_reg, col_reg}<14'b00001110111100)) color_data = 12'b010000100011;
		if(({row_reg, col_reg}==14'b00001110111100)) color_data = 12'b001100010100;
		if(({row_reg, col_reg}==14'b00001110111101)) color_data = 12'b001000000101;
		if(({row_reg, col_reg}==14'b00001110111110)) color_data = 12'b000100000111;
		if(({row_reg, col_reg}==14'b00001110111111)) color_data = 12'b000000001001;
		if(({row_reg, col_reg}>=14'b00001111000000) && ({row_reg, col_reg}<14'b00001111000011)) color_data = 12'b000000001110;

		if(({row_reg, col_reg}>=14'b00001111000011) && ({row_reg, col_reg}<14'b00010000101110)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=14'b00010000101110) && ({row_reg, col_reg}<14'b00010000110000)) color_data = 12'b000000001110;
		if(({row_reg, col_reg}==14'b00010000110000)) color_data = 12'b000100000101;
		if(({row_reg, col_reg}==14'b00010000110001)) color_data = 12'b001100100101;
		if(({row_reg, col_reg}==14'b00010000110010)) color_data = 12'b010100110100;
		if(({row_reg, col_reg}==14'b00010000110011)) color_data = 12'b010100100011;
		if(({row_reg, col_reg}==14'b00010000110100)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}==14'b00010000110101)) color_data = 12'b010100100011;
		if(({row_reg, col_reg}>=14'b00010000110110) && ({row_reg, col_reg}<14'b00010000111001)) color_data = 12'b010000100011;
		if(({row_reg, col_reg}>=14'b00010000111001) && ({row_reg, col_reg}<14'b00010000111100)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}==14'b00010000111100)) color_data = 12'b010000100011;
		if(({row_reg, col_reg}==14'b00010000111101)) color_data = 12'b001100100100;
		if(({row_reg, col_reg}==14'b00010000111110)) color_data = 12'b001000000101;
		if(({row_reg, col_reg}==14'b00010000111111)) color_data = 12'b000000000110;
		if(({row_reg, col_reg}>=14'b00010001000000) && ({row_reg, col_reg}<14'b00010001000010)) color_data = 12'b000000001100;
		if(({row_reg, col_reg}>=14'b00010001000010) && ({row_reg, col_reg}<14'b00010001000100)) color_data = 12'b000000001101;
		if(({row_reg, col_reg}==14'b00010001000100)) color_data = 12'b000000001110;

		if(({row_reg, col_reg}>=14'b00010001000101) && ({row_reg, col_reg}<14'b00010010101110)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=14'b00010010101110) && ({row_reg, col_reg}<14'b00010010110000)) color_data = 12'b000000001110;
		if(({row_reg, col_reg}==14'b00010010110000)) color_data = 12'b000100000110;
		if(({row_reg, col_reg}==14'b00010010110001)) color_data = 12'b001100100110;
		if(({row_reg, col_reg}==14'b00010010110010)) color_data = 12'b010100110101;
		if(({row_reg, col_reg}==14'b00010010110011)) color_data = 12'b010100100011;
		if(({row_reg, col_reg}==14'b00010010110100)) color_data = 12'b010100100010;
		if(({row_reg, col_reg}==14'b00010010110101)) color_data = 12'b010100100011;
		if(({row_reg, col_reg}>=14'b00010010110110) && ({row_reg, col_reg}<14'b00010010111010)) color_data = 12'b010000100011;
		if(({row_reg, col_reg}>=14'b00010010111010) && ({row_reg, col_reg}<14'b00010010111101)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}==14'b00010010111101)) color_data = 12'b010000100011;
		if(({row_reg, col_reg}==14'b00010010111110)) color_data = 12'b001100010100;
		if(({row_reg, col_reg}==14'b00010010111111)) color_data = 12'b001000000101;
		if(({row_reg, col_reg}==14'b00010011000000)) color_data = 12'b000100001000;
		if(({row_reg, col_reg}==14'b00010011000001)) color_data = 12'b000000001000;
		if(({row_reg, col_reg}==14'b00010011000010)) color_data = 12'b000000001001;
		if(({row_reg, col_reg}==14'b00010011000011)) color_data = 12'b000000001011;
		if(({row_reg, col_reg}==14'b00010011000100)) color_data = 12'b000000001100;
		if(({row_reg, col_reg}>=14'b00010011000101) && ({row_reg, col_reg}<14'b00010011000111)) color_data = 12'b000000001110;

		if(({row_reg, col_reg}>=14'b00010011000111) && ({row_reg, col_reg}<14'b00010100101110)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=14'b00010100101110) && ({row_reg, col_reg}<14'b00010100110000)) color_data = 12'b000000001110;
		if(({row_reg, col_reg}==14'b00010100110000)) color_data = 12'b000000000111;
		if(({row_reg, col_reg}==14'b00010100110001)) color_data = 12'b001000010110;
		if(({row_reg, col_reg}==14'b00010100110010)) color_data = 12'b001100100101;
		if(({row_reg, col_reg}==14'b00010100110011)) color_data = 12'b010000100100;
		if(({row_reg, col_reg}==14'b00010100110100)) color_data = 12'b010100100011;
		if(({row_reg, col_reg}>=14'b00010100110101) && ({row_reg, col_reg}<14'b00010100110111)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}>=14'b00010100110111) && ({row_reg, col_reg}<14'b00010100111011)) color_data = 12'b010000100011;
		if(({row_reg, col_reg}>=14'b00010100111011) && ({row_reg, col_reg}<14'b00010100111101)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}>=14'b00010100111101) && ({row_reg, col_reg}<14'b00010100111111)) color_data = 12'b010000100011;
		if(({row_reg, col_reg}==14'b00010100111111)) color_data = 12'b001100100100;
		if(({row_reg, col_reg}>=14'b00010101000000) && ({row_reg, col_reg}<14'b00010101000010)) color_data = 12'b000100000101;
		if(({row_reg, col_reg}==14'b00010101000010)) color_data = 12'b000100000110;
		if(({row_reg, col_reg}==14'b00010101000011)) color_data = 12'b000000000111;
		if(({row_reg, col_reg}==14'b00010101000100)) color_data = 12'b000000001001;
		if(({row_reg, col_reg}==14'b00010101000101)) color_data = 12'b000000001011;
		if(({row_reg, col_reg}==14'b00010101000110)) color_data = 12'b000000001101;
		if(({row_reg, col_reg}>=14'b00010101000111) && ({row_reg, col_reg}<14'b00010101001001)) color_data = 12'b000000001110;

		if(({row_reg, col_reg}>=14'b00010101001001) && ({row_reg, col_reg}<14'b00010110101111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==14'b00010110101111)) color_data = 12'b000000001110;
		if(({row_reg, col_reg}==14'b00010110110000)) color_data = 12'b000000001001;
		if(({row_reg, col_reg}==14'b00010110110001)) color_data = 12'b000100001000;
		if(({row_reg, col_reg}==14'b00010110110010)) color_data = 12'b001000010110;
		if(({row_reg, col_reg}==14'b00010110110011)) color_data = 12'b010000100101;
		if(({row_reg, col_reg}==14'b00010110110100)) color_data = 12'b010100110100;
		if(({row_reg, col_reg}==14'b00010110110101)) color_data = 12'b010100100011;
		if(({row_reg, col_reg}==14'b00010110110110)) color_data = 12'b010100100010;
		if(({row_reg, col_reg}==14'b00010110110111)) color_data = 12'b010100110011;
		if(({row_reg, col_reg}==14'b00010110111000)) color_data = 12'b010000100011;
		if(({row_reg, col_reg}>=14'b00010110111001) && ({row_reg, col_reg}<14'b00010110111011)) color_data = 12'b010000100100;
		if(({row_reg, col_reg}==14'b00010110111011)) color_data = 12'b010000100011;
		if(({row_reg, col_reg}>=14'b00010110111100) && ({row_reg, col_reg}<14'b00010110111111)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}==14'b00010110111111)) color_data = 12'b001100100011;
		if(({row_reg, col_reg}==14'b00010111000000)) color_data = 12'b010000100011;
		if(({row_reg, col_reg}==14'b00010111000001)) color_data = 12'b010000100100;
		if(({row_reg, col_reg}==14'b00010111000010)) color_data = 12'b001100010101;
		if(({row_reg, col_reg}==14'b00010111000011)) color_data = 12'b001000010101;
		if(({row_reg, col_reg}==14'b00010111000100)) color_data = 12'b000100000111;
		if(({row_reg, col_reg}==14'b00010111000101)) color_data = 12'b000000001000;
		if(({row_reg, col_reg}==14'b00010111000110)) color_data = 12'b000000001010;
		if(({row_reg, col_reg}>=14'b00010111000111) && ({row_reg, col_reg}<14'b00010111001001)) color_data = 12'b000000001100;
		if(({row_reg, col_reg}==14'b00010111001001)) color_data = 12'b000000001110;

		if(({row_reg, col_reg}>=14'b00010111001010) && ({row_reg, col_reg}<14'b00011000110000)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==14'b00011000110000)) color_data = 12'b000000001100;
		if(({row_reg, col_reg}==14'b00011000110001)) color_data = 12'b000000001010;
		if(({row_reg, col_reg}==14'b00011000110010)) color_data = 12'b000100001000;
		if(({row_reg, col_reg}==14'b00011000110011)) color_data = 12'b001000010110;
		if(({row_reg, col_reg}==14'b00011000110100)) color_data = 12'b010000100101;
		if(({row_reg, col_reg}==14'b00011000110101)) color_data = 12'b010100100100;
		if(({row_reg, col_reg}==14'b00011000110110)) color_data = 12'b010100100011;
		if(({row_reg, col_reg}>=14'b00011000110111) && ({row_reg, col_reg}<14'b00011000111001)) color_data = 12'b010000100011;
		if(({row_reg, col_reg}>=14'b00011000111001) && ({row_reg, col_reg}<14'b00011000111011)) color_data = 12'b010000100100;
		if(({row_reg, col_reg}>=14'b00011000111011) && ({row_reg, col_reg}<14'b00011000111101)) color_data = 12'b010000100011;
		if(({row_reg, col_reg}>=14'b00011000111101) && ({row_reg, col_reg}<14'b00011001000010)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}==14'b00011001000010)) color_data = 12'b010000100011;
		if(({row_reg, col_reg}==14'b00011001000011)) color_data = 12'b001100010100;
		if(({row_reg, col_reg}==14'b00011001000100)) color_data = 12'b001000010101;
		if(({row_reg, col_reg}==14'b00011001000101)) color_data = 12'b000100000101;
		if(({row_reg, col_reg}==14'b00011001000110)) color_data = 12'b000100000110;
		if(({row_reg, col_reg}==14'b00011001000111)) color_data = 12'b000000001000;
		if(({row_reg, col_reg}==14'b00011001001000)) color_data = 12'b000000001001;
		if(({row_reg, col_reg}==14'b00011001001001)) color_data = 12'b000000001011;
		if(({row_reg, col_reg}==14'b00011001001010)) color_data = 12'b000000001101;
		if(({row_reg, col_reg}==14'b00011001001011)) color_data = 12'b000000001110;

		if(({row_reg, col_reg}>=14'b00011001001100) && ({row_reg, col_reg}<14'b00011010110000)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==14'b00011010110000)) color_data = 12'b000000001110;
		if(({row_reg, col_reg}==14'b00011010110001)) color_data = 12'b000000001101;
		if(({row_reg, col_reg}==14'b00011010110010)) color_data = 12'b000000001010;
		if(({row_reg, col_reg}==14'b00011010110011)) color_data = 12'b000000000111;
		if(({row_reg, col_reg}==14'b00011010110100)) color_data = 12'b001000000110;
		if(({row_reg, col_reg}==14'b00011010110101)) color_data = 12'b001100100110;
		if(({row_reg, col_reg}==14'b00011010110110)) color_data = 12'b010000100100;
		if(({row_reg, col_reg}>=14'b00011010110111) && ({row_reg, col_reg}<14'b00011010111010)) color_data = 12'b010000100011;
		if(({row_reg, col_reg}==14'b00011010111010)) color_data = 12'b010000100100;
		if(({row_reg, col_reg}>=14'b00011010111011) && ({row_reg, col_reg}<14'b00011010111101)) color_data = 12'b010000100011;
		if(({row_reg, col_reg}>=14'b00011010111101) && ({row_reg, col_reg}<14'b00011011000011)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}==14'b00011011000011)) color_data = 12'b010000100011;
		if(({row_reg, col_reg}==14'b00011011000100)) color_data = 12'b010000100100;
		if(({row_reg, col_reg}==14'b00011011000101)) color_data = 12'b001100100100;
		if(({row_reg, col_reg}==14'b00011011000110)) color_data = 12'b001100010101;
		if(({row_reg, col_reg}==14'b00011011000111)) color_data = 12'b001000010110;
		if(({row_reg, col_reg}==14'b00011011001000)) color_data = 12'b000000000110;
		if(({row_reg, col_reg}==14'b00011011001001)) color_data = 12'b000000001000;
		if(({row_reg, col_reg}==14'b00011011001010)) color_data = 12'b000000001010;
		if(({row_reg, col_reg}==14'b00011011001011)) color_data = 12'b000000001100;
		if(({row_reg, col_reg}==14'b00011011001100)) color_data = 12'b000000001110;

		if(({row_reg, col_reg}>=14'b00011011001101) && ({row_reg, col_reg}<14'b00011100110010)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==14'b00011100110010)) color_data = 12'b000000001101;
		if(({row_reg, col_reg}==14'b00011100110011)) color_data = 12'b000000001011;
		if(({row_reg, col_reg}==14'b00011100110100)) color_data = 12'b000100001001;
		if(({row_reg, col_reg}==14'b00011100110101)) color_data = 12'b001000000111;
		if(({row_reg, col_reg}==14'b00011100110110)) color_data = 12'b001100100101;
		if(({row_reg, col_reg}==14'b00011100110111)) color_data = 12'b010000100100;
		if(({row_reg, col_reg}==14'b00011100111000)) color_data = 12'b010000100011;
		if(({row_reg, col_reg}==14'b00011100111001)) color_data = 12'b010100100011;
		if(({row_reg, col_reg}>=14'b00011100111010) && ({row_reg, col_reg}<14'b00011101000010)) color_data = 12'b010000100011;
		if(({row_reg, col_reg}==14'b00011101000010)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}==14'b00011101000011)) color_data = 12'b010000010010;
		if(({row_reg, col_reg}==14'b00011101000100)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}>=14'b00011101000101) && ({row_reg, col_reg}<14'b00011101000111)) color_data = 12'b010000100011;
		if(({row_reg, col_reg}==14'b00011101000111)) color_data = 12'b001100100011;
		if(({row_reg, col_reg}==14'b00011101001000)) color_data = 12'b001000010100;
		if(({row_reg, col_reg}==14'b00011101001001)) color_data = 12'b000100000101;
		if(({row_reg, col_reg}==14'b00011101001010)) color_data = 12'b000100001000;
		if(({row_reg, col_reg}==14'b00011101001011)) color_data = 12'b000000001010;
		if(({row_reg, col_reg}==14'b00011101001100)) color_data = 12'b000000001101;

		if(({row_reg, col_reg}>=14'b00011101001101) && ({row_reg, col_reg}<14'b00011110110010)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==14'b00011110110010)) color_data = 12'b000000001110;
		if(({row_reg, col_reg}==14'b00011110110011)) color_data = 12'b000100001101;
		if(({row_reg, col_reg}==14'b00011110110100)) color_data = 12'b000100001010;
		if(({row_reg, col_reg}==14'b00011110110101)) color_data = 12'b000000000111;
		if(({row_reg, col_reg}==14'b00011110110110)) color_data = 12'b000100000101;
		if(({row_reg, col_reg}==14'b00011110110111)) color_data = 12'b010000100101;
		if(({row_reg, col_reg}==14'b00011110111000)) color_data = 12'b010000100011;
		if(({row_reg, col_reg}>=14'b00011110111001) && ({row_reg, col_reg}<14'b00011110111100)) color_data = 12'b010100100011;
		if(({row_reg, col_reg}>=14'b00011110111100) && ({row_reg, col_reg}<14'b00011111000000)) color_data = 12'b010000100011;
		if(({row_reg, col_reg}==14'b00011111000000)) color_data = 12'b010000100100;
		if(({row_reg, col_reg}>=14'b00011111000001) && ({row_reg, col_reg}<14'b00011111000011)) color_data = 12'b010000100011;
		if(({row_reg, col_reg}>=14'b00011111000011) && ({row_reg, col_reg}<14'b00011111000110)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}==14'b00011111000110)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==14'b00011111000111)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}==14'b00011111001000)) color_data = 12'b010000100011;
		if(({row_reg, col_reg}==14'b00011111001001)) color_data = 12'b001100010100;
		if(({row_reg, col_reg}==14'b00011111001010)) color_data = 12'b000100000110;
		if(({row_reg, col_reg}==14'b00011111001011)) color_data = 12'b000000001001;
		if(({row_reg, col_reg}==14'b00011111001100)) color_data = 12'b000000001100;
		if(({row_reg, col_reg}==14'b00011111001101)) color_data = 12'b000000001110;

		if(({row_reg, col_reg}>=14'b00011111001110) && ({row_reg, col_reg}<14'b00100000110100)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==14'b00100000110100)) color_data = 12'b000000001110;
		if(({row_reg, col_reg}==14'b00100000110101)) color_data = 12'b000000001100;
		if(({row_reg, col_reg}==14'b00100000110110)) color_data = 12'b000100001001;
		if(({row_reg, col_reg}==14'b00100000110111)) color_data = 12'b000100000110;
		if(({row_reg, col_reg}==14'b00100000111000)) color_data = 12'b010000100110;
		if(({row_reg, col_reg}==14'b00100000111001)) color_data = 12'b010000100100;
		if(({row_reg, col_reg}>=14'b00100000111010) && ({row_reg, col_reg}<14'b00100000111101)) color_data = 12'b010100100011;
		if(({row_reg, col_reg}>=14'b00100000111101) && ({row_reg, col_reg}<14'b00100000111111)) color_data = 12'b010000100011;
		if(({row_reg, col_reg}==14'b00100000111111)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}==14'b00100001000000)) color_data = 12'b010000100011;
		if(({row_reg, col_reg}>=14'b00100001000001) && ({row_reg, col_reg}<14'b00100001000011)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}>=14'b00100001000011) && ({row_reg, col_reg}<14'b00100001000101)) color_data = 12'b010000100011;
		if(({row_reg, col_reg}>=14'b00100001000101) && ({row_reg, col_reg}<14'b00100001000111)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}>=14'b00100001000111) && ({row_reg, col_reg}<14'b00100001001001)) color_data = 12'b010000100011;
		if(({row_reg, col_reg}==14'b00100001001001)) color_data = 12'b001100010011;
		if(({row_reg, col_reg}==14'b00100001001010)) color_data = 12'b001000010011;
		if(({row_reg, col_reg}==14'b00100001001011)) color_data = 12'b001000000101;
		if(({row_reg, col_reg}==14'b00100001001100)) color_data = 12'b000100000111;
		if(({row_reg, col_reg}==14'b00100001001101)) color_data = 12'b000000001010;
		if(({row_reg, col_reg}==14'b00100001001110)) color_data = 12'b000000001110;

		if(({row_reg, col_reg}>=14'b00100001001111) && ({row_reg, col_reg}<14'b00100010110101)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==14'b00100010110101)) color_data = 12'b000000001101;
		if(({row_reg, col_reg}==14'b00100010110110)) color_data = 12'b000000001011;
		if(({row_reg, col_reg}==14'b00100010110111)) color_data = 12'b000100001000;
		if(({row_reg, col_reg}==14'b00100010111000)) color_data = 12'b001000000101;
		if(({row_reg, col_reg}==14'b00100010111001)) color_data = 12'b001100010100;
		if(({row_reg, col_reg}==14'b00100010111010)) color_data = 12'b010100100100;
		if(({row_reg, col_reg}==14'b00100010111011)) color_data = 12'b010100100011;
		if(({row_reg, col_reg}>=14'b00100010111100) && ({row_reg, col_reg}<14'b00100010111110)) color_data = 12'b010000100011;
		if(({row_reg, col_reg}==14'b00100010111110)) color_data = 12'b010100100011;
		if(({row_reg, col_reg}==14'b00100010111111)) color_data = 12'b010000100011;
		if(({row_reg, col_reg}>=14'b00100011000000) && ({row_reg, col_reg}<14'b00100011000011)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}>=14'b00100011000011) && ({row_reg, col_reg}<14'b00100011000110)) color_data = 12'b010000100011;
		if(({row_reg, col_reg}>=14'b00100011000110) && ({row_reg, col_reg}<14'b00100011001001)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}==14'b00100011001001)) color_data = 12'b010000100011;
		if(({row_reg, col_reg}==14'b00100011001010)) color_data = 12'b010000100100;
		if(({row_reg, col_reg}==14'b00100011001011)) color_data = 12'b001100010100;
		if(({row_reg, col_reg}==14'b00100011001100)) color_data = 12'b000100000110;
		if(({row_reg, col_reg}==14'b00100011001101)) color_data = 12'b000000001000;
		if(({row_reg, col_reg}==14'b00100011001110)) color_data = 12'b000000001011;
		if(({row_reg, col_reg}>=14'b00100011001111) && ({row_reg, col_reg}<14'b00100011010001)) color_data = 12'b000000001110;

		if(({row_reg, col_reg}>=14'b00100011010001) && ({row_reg, col_reg}<14'b00100100110101)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==14'b00100100110101)) color_data = 12'b000000001110;
		if(({row_reg, col_reg}==14'b00100100110110)) color_data = 12'b000000001101;
		if(({row_reg, col_reg}==14'b00100100110111)) color_data = 12'b000100001010;
		if(({row_reg, col_reg}==14'b00100100111000)) color_data = 12'b000100000111;
		if(({row_reg, col_reg}==14'b00100100111001)) color_data = 12'b001000010110;
		if(({row_reg, col_reg}==14'b00100100111010)) color_data = 12'b010000100101;
		if(({row_reg, col_reg}==14'b00100100111011)) color_data = 12'b010000100100;
		if(({row_reg, col_reg}>=14'b00100100111100) && ({row_reg, col_reg}<14'b00100101000110)) color_data = 12'b010000100011;
		if(({row_reg, col_reg}>=14'b00100101000110) && ({row_reg, col_reg}<14'b00100101001000)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}==14'b00100101001000)) color_data = 12'b010000010010;
		if(({row_reg, col_reg}==14'b00100101001001)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}==14'b00100101001010)) color_data = 12'b010000100011;
		if(({row_reg, col_reg}==14'b00100101001011)) color_data = 12'b010000010011;
		if(({row_reg, col_reg}==14'b00100101001100)) color_data = 12'b001100010100;
		if(({row_reg, col_reg}==14'b00100101001101)) color_data = 12'b001000000110;
		if(({row_reg, col_reg}==14'b00100101001110)) color_data = 12'b000100001000;
		if(({row_reg, col_reg}==14'b00100101001111)) color_data = 12'b000000001001;
		if(({row_reg, col_reg}==14'b00100101010000)) color_data = 12'b000000001010;
		if(({row_reg, col_reg}==14'b00100101010001)) color_data = 12'b000000001011;
		if(({row_reg, col_reg}==14'b00100101010010)) color_data = 12'b000000001101;

		if(({row_reg, col_reg}>=14'b00100101010011) && ({row_reg, col_reg}<14'b00100110110110)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==14'b00100110110110)) color_data = 12'b000000001110;
		if(({row_reg, col_reg}==14'b00100110110111)) color_data = 12'b000000001101;
		if(({row_reg, col_reg}==14'b00100110111000)) color_data = 12'b000100001010;
		if(({row_reg, col_reg}==14'b00100110111001)) color_data = 12'b000100001000;
		if(({row_reg, col_reg}==14'b00100110111010)) color_data = 12'b001000010110;
		if(({row_reg, col_reg}==14'b00100110111011)) color_data = 12'b001100100101;
		if(({row_reg, col_reg}>=14'b00100110111100) && ({row_reg, col_reg}<14'b00100110111110)) color_data = 12'b010000100100;
		if(({row_reg, col_reg}==14'b00100110111110)) color_data = 12'b010000100011;
		if(({row_reg, col_reg}==14'b00100110111111)) color_data = 12'b010100100011;
		if(({row_reg, col_reg}==14'b00100111000000)) color_data = 12'b010000100011;
		if(({row_reg, col_reg}>=14'b00100111000001) && ({row_reg, col_reg}<14'b00100111000011)) color_data = 12'b010100100011;
		if(({row_reg, col_reg}>=14'b00100111000011) && ({row_reg, col_reg}<14'b00100111000111)) color_data = 12'b010000100011;
		if(({row_reg, col_reg}>=14'b00100111000111) && ({row_reg, col_reg}<14'b00100111001010)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}>=14'b00100111001010) && ({row_reg, col_reg}<14'b00100111001101)) color_data = 12'b010000100011;
		if(({row_reg, col_reg}==14'b00100111001101)) color_data = 12'b001100010100;
		if(({row_reg, col_reg}==14'b00100111001110)) color_data = 12'b001000000100;
		if(({row_reg, col_reg}==14'b00100111001111)) color_data = 12'b000100000101;
		if(({row_reg, col_reg}==14'b00100111010000)) color_data = 12'b000100000111;
		if(({row_reg, col_reg}==14'b00100111010001)) color_data = 12'b000000001000;
		if(({row_reg, col_reg}==14'b00100111010010)) color_data = 12'b000000001010;
		if(({row_reg, col_reg}==14'b00100111010011)) color_data = 12'b000000001101;

		if(({row_reg, col_reg}>=14'b00100111010100) && ({row_reg, col_reg}<14'b00101000111000)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==14'b00101000111000)) color_data = 12'b000000001101;
		if(({row_reg, col_reg}==14'b00101000111001)) color_data = 12'b000000001010;
		if(({row_reg, col_reg}==14'b00101000111010)) color_data = 12'b000100001000;
		if(({row_reg, col_reg}==14'b00101000111011)) color_data = 12'b001000010110;
		if(({row_reg, col_reg}==14'b00101000111100)) color_data = 12'b001100100101;
		if(({row_reg, col_reg}==14'b00101000111101)) color_data = 12'b010000100100;
		if(({row_reg, col_reg}==14'b00101000111110)) color_data = 12'b010100100100;
		if(({row_reg, col_reg}==14'b00101000111111)) color_data = 12'b010100100011;
		if(({row_reg, col_reg}>=14'b00101001000000) && ({row_reg, col_reg}<14'b00101001000111)) color_data = 12'b010000100011;
		if(({row_reg, col_reg}>=14'b00101001000111) && ({row_reg, col_reg}<14'b00101001001010)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}>=14'b00101001001010) && ({row_reg, col_reg}<14'b00101001001110)) color_data = 12'b010000100011;
		if(({row_reg, col_reg}>=14'b00101001001110) && ({row_reg, col_reg}<14'b00101001010000)) color_data = 12'b001100100100;
		if(({row_reg, col_reg}==14'b00101001010000)) color_data = 12'b001000010100;
		if(({row_reg, col_reg}==14'b00101001010001)) color_data = 12'b000100000101;
		if(({row_reg, col_reg}==14'b00101001010010)) color_data = 12'b000100000111;
		if(({row_reg, col_reg}==14'b00101001010011)) color_data = 12'b000000001011;
		if(({row_reg, col_reg}==14'b00101001010100)) color_data = 12'b000000001101;
		if(({row_reg, col_reg}==14'b00101001010101)) color_data = 12'b000000001110;

		if(({row_reg, col_reg}>=14'b00101001010110) && ({row_reg, col_reg}<14'b00101010111001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==14'b00101010111001)) color_data = 12'b000000001101;
		if(({row_reg, col_reg}==14'b00101010111010)) color_data = 12'b000000001011;
		if(({row_reg, col_reg}==14'b00101010111011)) color_data = 12'b000000001000;
		if(({row_reg, col_reg}==14'b00101010111100)) color_data = 12'b001000000110;
		if(({row_reg, col_reg}==14'b00101010111101)) color_data = 12'b001100100101;
		if(({row_reg, col_reg}==14'b00101010111110)) color_data = 12'b010000100100;
		if(({row_reg, col_reg}==14'b00101010111111)) color_data = 12'b010100100011;
		if(({row_reg, col_reg}==14'b00101011000000)) color_data = 12'b010000100011;
		if(({row_reg, col_reg}>=14'b00101011000001) && ({row_reg, col_reg}<14'b00101011000011)) color_data = 12'b010100100011;
		if(({row_reg, col_reg}==14'b00101011000011)) color_data = 12'b010100100100;
		if(({row_reg, col_reg}==14'b00101011000100)) color_data = 12'b010000100100;
		if(({row_reg, col_reg}>=14'b00101011000101) && ({row_reg, col_reg}<14'b00101011001100)) color_data = 12'b010000100011;
		if(({row_reg, col_reg}>=14'b00101011001100) && ({row_reg, col_reg}<14'b00101011001111)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}==14'b00101011001111)) color_data = 12'b010000100011;
		if(({row_reg, col_reg}==14'b00101011010000)) color_data = 12'b001100100011;
		if(({row_reg, col_reg}==14'b00101011010001)) color_data = 12'b001100010100;
		if(({row_reg, col_reg}==14'b00101011010010)) color_data = 12'b000100000101;
		if(({row_reg, col_reg}==14'b00101011010011)) color_data = 12'b000000000111;
		if(({row_reg, col_reg}==14'b00101011010100)) color_data = 12'b000000001010;
		if(({row_reg, col_reg}==14'b00101011010101)) color_data = 12'b000000001100;
		if(({row_reg, col_reg}==14'b00101011010110)) color_data = 12'b000000001110;

		if(({row_reg, col_reg}>=14'b00101011010111) && ({row_reg, col_reg}<14'b00101100111010)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==14'b00101100111010)) color_data = 12'b000000001101;
		if(({row_reg, col_reg}==14'b00101100111011)) color_data = 12'b000000001011;
		if(({row_reg, col_reg}==14'b00101100111100)) color_data = 12'b000100001000;
		if(({row_reg, col_reg}==14'b00101100111101)) color_data = 12'b001000000110;
		if(({row_reg, col_reg}==14'b00101100111110)) color_data = 12'b001100010100;
		if(({row_reg, col_reg}==14'b00101100111111)) color_data = 12'b010000100100;
		if(({row_reg, col_reg}==14'b00101101000000)) color_data = 12'b010100100100;
		if(({row_reg, col_reg}>=14'b00101101000001) && ({row_reg, col_reg}<14'b00101101000100)) color_data = 12'b010100100011;
		if(({row_reg, col_reg}>=14'b00101101000100) && ({row_reg, col_reg}<14'b00101101000110)) color_data = 12'b010000100011;
		if(({row_reg, col_reg}>=14'b00101101000110) && ({row_reg, col_reg}<14'b00101101001000)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}==14'b00101101001000)) color_data = 12'b010000010010;
		if(({row_reg, col_reg}==14'b00101101001001)) color_data = 12'b001100010010;
		if(({row_reg, col_reg}==14'b00101101001010)) color_data = 12'b001100100011;
		if(({row_reg, col_reg}>=14'b00101101001011) && ({row_reg, col_reg}<14'b00101101001101)) color_data = 12'b010000100011;
		if(({row_reg, col_reg}>=14'b00101101001101) && ({row_reg, col_reg}<14'b00101101010001)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}==14'b00101101010001)) color_data = 12'b001100100011;
		if(({row_reg, col_reg}==14'b00101101010010)) color_data = 12'b001100010100;
		if(({row_reg, col_reg}==14'b00101101010011)) color_data = 12'b000100000101;
		if(({row_reg, col_reg}==14'b00101101010100)) color_data = 12'b000000000111;
		if(({row_reg, col_reg}==14'b00101101010101)) color_data = 12'b000000001010;
		if(({row_reg, col_reg}==14'b00101101010110)) color_data = 12'b000000001100;
		if(({row_reg, col_reg}==14'b00101101010111)) color_data = 12'b000000001110;

		if(({row_reg, col_reg}>=14'b00101101011000) && ({row_reg, col_reg}<14'b00101110111011)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==14'b00101110111011)) color_data = 12'b000000001101;
		if(({row_reg, col_reg}==14'b00101110111100)) color_data = 12'b000000001011;
		if(({row_reg, col_reg}==14'b00101110111101)) color_data = 12'b000100001000;
		if(({row_reg, col_reg}==14'b00101110111110)) color_data = 12'b001000010110;
		if(({row_reg, col_reg}==14'b00101110111111)) color_data = 12'b010000100110;
		if(({row_reg, col_reg}==14'b00101111000000)) color_data = 12'b010000100100;
		if(({row_reg, col_reg}==14'b00101111000001)) color_data = 12'b010000100011;
		if(({row_reg, col_reg}==14'b00101111000010)) color_data = 12'b010000010010;
		if(({row_reg, col_reg}>=14'b00101111000011) && ({row_reg, col_reg}<14'b00101111000101)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}==14'b00101111000101)) color_data = 12'b001100010010;
		if(({row_reg, col_reg}>=14'b00101111000110) && ({row_reg, col_reg}<14'b00101111001001)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}==14'b00101111001001)) color_data = 12'b010000100011;
		if(({row_reg, col_reg}==14'b00101111001010)) color_data = 12'b001100100011;
		if(({row_reg, col_reg}>=14'b00101111001011) && ({row_reg, col_reg}<14'b00101111001101)) color_data = 12'b010000100011;
		if(({row_reg, col_reg}>=14'b00101111001101) && ({row_reg, col_reg}<14'b00101111010010)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}==14'b00101111010010)) color_data = 12'b010000100011;
		if(({row_reg, col_reg}==14'b00101111010011)) color_data = 12'b001100010100;
		if(({row_reg, col_reg}==14'b00101111010100)) color_data = 12'b000100010101;
		if(({row_reg, col_reg}==14'b00101111010101)) color_data = 12'b000100001000;
		if(({row_reg, col_reg}==14'b00101111010110)) color_data = 12'b000000001010;
		if(({row_reg, col_reg}==14'b00101111010111)) color_data = 12'b000000001101;

		if(({row_reg, col_reg}>=14'b00101111011000) && ({row_reg, col_reg}<14'b00110000111100)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==14'b00110000111100)) color_data = 12'b000000001101;
		if(({row_reg, col_reg}==14'b00110000111101)) color_data = 12'b000000001010;
		if(({row_reg, col_reg}==14'b00110000111110)) color_data = 12'b000100001000;
		if(({row_reg, col_reg}==14'b00110000111111)) color_data = 12'b000100000110;
		if(({row_reg, col_reg}==14'b00110001000000)) color_data = 12'b001100010100;
		if(({row_reg, col_reg}==14'b00110001000001)) color_data = 12'b001100010011;
		if(({row_reg, col_reg}==14'b00110001000010)) color_data = 12'b001100010010;
		if(({row_reg, col_reg}>=14'b00110001000011) && ({row_reg, col_reg}<14'b00110001000101)) color_data = 12'b001100010001;
		if(({row_reg, col_reg}>=14'b00110001000101) && ({row_reg, col_reg}<14'b00110001000111)) color_data = 12'b001100010010;
		if(({row_reg, col_reg}>=14'b00110001000111) && ({row_reg, col_reg}<14'b00110001001001)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}==14'b00110001001001)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}>=14'b00110001001010) && ({row_reg, col_reg}<14'b00110001001100)) color_data = 12'b001100100011;
		if(({row_reg, col_reg}==14'b00110001001100)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==14'b00110001001101)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}==14'b00110001001110)) color_data = 12'b010000100011;
		if(({row_reg, col_reg}==14'b00110001001111)) color_data = 12'b010000010010;
		if(({row_reg, col_reg}>=14'b00110001010000) && ({row_reg, col_reg}<14'b00110001010011)) color_data = 12'b010000100011;
		if(({row_reg, col_reg}==14'b00110001010011)) color_data = 12'b001100100011;
		if(({row_reg, col_reg}==14'b00110001010100)) color_data = 12'b001100100100;
		if(({row_reg, col_reg}==14'b00110001010101)) color_data = 12'b000100000101;
		if(({row_reg, col_reg}==14'b00110001010110)) color_data = 12'b000000000111;
		if(({row_reg, col_reg}==14'b00110001010111)) color_data = 12'b000100001011;
		if(({row_reg, col_reg}==14'b00110001011000)) color_data = 12'b000000001110;

		if(({row_reg, col_reg}>=14'b00110001011001) && ({row_reg, col_reg}<14'b00110010111100)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==14'b00110010111100)) color_data = 12'b000000001110;
		if(({row_reg, col_reg}==14'b00110010111101)) color_data = 12'b000000001100;
		if(({row_reg, col_reg}==14'b00110010111110)) color_data = 12'b000000001010;
		if(({row_reg, col_reg}==14'b00110010111111)) color_data = 12'b000000001001;
		if(({row_reg, col_reg}==14'b00110011000000)) color_data = 12'b001000000100;
		if(({row_reg, col_reg}==14'b00110011000001)) color_data = 12'b001100010100;
		if(({row_reg, col_reg}==14'b00110011000010)) color_data = 12'b010100100100;
		if(({row_reg, col_reg}==14'b00110011000011)) color_data = 12'b011000110100;
		if(({row_reg, col_reg}==14'b00110011000100)) color_data = 12'b010100110011;
		if(({row_reg, col_reg}==14'b00110011000101)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==14'b00110011000110)) color_data = 12'b001100010010;
		if(({row_reg, col_reg}==14'b00110011000111)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}>=14'b00110011001000) && ({row_reg, col_reg}<14'b00110011001010)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}>=14'b00110011001010) && ({row_reg, col_reg}<14'b00110011001100)) color_data = 12'b001100100011;
		if(({row_reg, col_reg}>=14'b00110011001100) && ({row_reg, col_reg}<14'b00110011010010)) color_data = 12'b010000100011;
		if(({row_reg, col_reg}==14'b00110011010010)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}==14'b00110011010011)) color_data = 12'b010000100011;
		if(({row_reg, col_reg}==14'b00110011010100)) color_data = 12'b010000100100;
		if(({row_reg, col_reg}==14'b00110011010101)) color_data = 12'b001100010100;
		if(({row_reg, col_reg}==14'b00110011010110)) color_data = 12'b000100000101;
		if(({row_reg, col_reg}==14'b00110011010111)) color_data = 12'b000100001000;
		if(({row_reg, col_reg}==14'b00110011011000)) color_data = 12'b000000001011;
		if(({row_reg, col_reg}==14'b00110011011001)) color_data = 12'b000000001101;

		if(({row_reg, col_reg}>=14'b00110011011010) && ({row_reg, col_reg}<14'b00110100111101)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==14'b00110100111101)) color_data = 12'b000000001110;
		if(({row_reg, col_reg}==14'b00110100111110)) color_data = 12'b000000001100;
		if(({row_reg, col_reg}==14'b00110100111111)) color_data = 12'b000000001011;
		if(({row_reg, col_reg}==14'b00110101000000)) color_data = 12'b000100000100;
		if(({row_reg, col_reg}==14'b00110101000001)) color_data = 12'b001000000011;
		if(({row_reg, col_reg}==14'b00110101000010)) color_data = 12'b011101000110;
		if(({row_reg, col_reg}==14'b00110101000011)) color_data = 12'b101001111000;
		if(({row_reg, col_reg}==14'b00110101000100)) color_data = 12'b100001010101;
		if(({row_reg, col_reg}==14'b00110101000101)) color_data = 12'b001100010010;
		if(({row_reg, col_reg}==14'b00110101000110)) color_data = 12'b001100010001;
		if(({row_reg, col_reg}==14'b00110101000111)) color_data = 12'b010000100011;
		if(({row_reg, col_reg}==14'b00110101001000)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}>=14'b00110101001001) && ({row_reg, col_reg}<14'b00110101001011)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}>=14'b00110101001011) && ({row_reg, col_reg}<14'b00110101001101)) color_data = 12'b001100100011;
		if(({row_reg, col_reg}>=14'b00110101001101) && ({row_reg, col_reg}<14'b00110101010110)) color_data = 12'b010000100011;
		if(({row_reg, col_reg}==14'b00110101010110)) color_data = 12'b001100010100;
		if(({row_reg, col_reg}==14'b00110101010111)) color_data = 12'b000100000101;
		if(({row_reg, col_reg}==14'b00110101011000)) color_data = 12'b000000000111;
		if(({row_reg, col_reg}==14'b00110101011001)) color_data = 12'b000000001010;
		if(({row_reg, col_reg}==14'b00110101011010)) color_data = 12'b000000001101;

		if(({row_reg, col_reg}>=14'b00110101011011) && ({row_reg, col_reg}<14'b00110110111110)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=14'b00110110111110) && ({row_reg, col_reg}<14'b00110111000000)) color_data = 12'b000000001101;
		if(({row_reg, col_reg}==14'b00110111000000)) color_data = 12'b001000000100;
		if(({row_reg, col_reg}==14'b00110111000001)) color_data = 12'b001100000011;
		if(({row_reg, col_reg}==14'b00110111000010)) color_data = 12'b100001000101;
		if(({row_reg, col_reg}==14'b00110111000011)) color_data = 12'b101001110111;
		if(({row_reg, col_reg}==14'b00110111000100)) color_data = 12'b100001000101;
		if(({row_reg, col_reg}==14'b00110111000101)) color_data = 12'b010100100011;
		if(({row_reg, col_reg}==14'b00110111000110)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}==14'b00110111000111)) color_data = 12'b001100010010;
		if(({row_reg, col_reg}==14'b00110111001000)) color_data = 12'b010000010010;
		if(({row_reg, col_reg}>=14'b00110111001001) && ({row_reg, col_reg}<14'b00110111001100)) color_data = 12'b001100010010;
		if(({row_reg, col_reg}==14'b00110111001100)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}>=14'b00110111001101) && ({row_reg, col_reg}<14'b00110111010000)) color_data = 12'b010000100011;
		if(({row_reg, col_reg}>=14'b00110111010000) && ({row_reg, col_reg}<14'b00110111010010)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}>=14'b00110111010010) && ({row_reg, col_reg}<14'b00110111010100)) color_data = 12'b010000100011;
		if(({row_reg, col_reg}==14'b00110111010100)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}>=14'b00110111010101) && ({row_reg, col_reg}<14'b00110111010111)) color_data = 12'b010000100011;
		if(({row_reg, col_reg}==14'b00110111010111)) color_data = 12'b001100010100;
		if(({row_reg, col_reg}==14'b00110111011000)) color_data = 12'b000100000101;
		if(({row_reg, col_reg}==14'b00110111011001)) color_data = 12'b000100001000;
		if(({row_reg, col_reg}==14'b00110111011010)) color_data = 12'b000000001011;
		if(({row_reg, col_reg}==14'b00110111011011)) color_data = 12'b000000001101;

		if(({row_reg, col_reg}>=14'b00110111011100) && ({row_reg, col_reg}<14'b00111000111110)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==14'b00111000111110)) color_data = 12'b000000001110;
		if(({row_reg, col_reg}==14'b00111000111111)) color_data = 12'b000000001101;
		if(({row_reg, col_reg}==14'b00111001000000)) color_data = 12'b001000000100;
		if(({row_reg, col_reg}==14'b00111001000001)) color_data = 12'b010000000011;
		if(({row_reg, col_reg}==14'b00111001000010)) color_data = 12'b011100100011;
		if(({row_reg, col_reg}>=14'b00111001000011) && ({row_reg, col_reg}<14'b00111001000101)) color_data = 12'b100000110011;
		if(({row_reg, col_reg}==14'b00111001000101)) color_data = 12'b100101100110;
		if(({row_reg, col_reg}==14'b00111001000110)) color_data = 12'b100101100111;
		if(({row_reg, col_reg}==14'b00111001000111)) color_data = 12'b010000100011;
		if(({row_reg, col_reg}==14'b00111001001000)) color_data = 12'b010000010010;
		if(({row_reg, col_reg}>=14'b00111001001001) && ({row_reg, col_reg}<14'b00111001001011)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}==14'b00111001001011)) color_data = 12'b001100010010;
		if(({row_reg, col_reg}>=14'b00111001001100) && ({row_reg, col_reg}<14'b00111001001110)) color_data = 12'b010000100011;
		if(({row_reg, col_reg}>=14'b00111001001110) && ({row_reg, col_reg}<14'b00111001010001)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}==14'b00111001010001)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}>=14'b00111001010010) && ({row_reg, col_reg}<14'b00111001010100)) color_data = 12'b010000100011;
		if(({row_reg, col_reg}>=14'b00111001010100) && ({row_reg, col_reg}<14'b00111001010111)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}==14'b00111001010111)) color_data = 12'b010000100011;
		if(({row_reg, col_reg}==14'b00111001011000)) color_data = 12'b001000010100;
		if(({row_reg, col_reg}==14'b00111001011001)) color_data = 12'b001000000110;
		if(({row_reg, col_reg}==14'b00111001011010)) color_data = 12'b000100001000;
		if(({row_reg, col_reg}==14'b00111001011011)) color_data = 12'b000000001010;
		if(({row_reg, col_reg}==14'b00111001011100)) color_data = 12'b000000001101;
		if(({row_reg, col_reg}==14'b00111001011101)) color_data = 12'b000000001110;

		if(({row_reg, col_reg}>=14'b00111001011110) && ({row_reg, col_reg}<14'b00111010111101)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==14'b00111010111101)) color_data = 12'b000000001110;
		if(({row_reg, col_reg}>=14'b00111010111110) && ({row_reg, col_reg}<14'b00111011000000)) color_data = 12'b000000001101;
		if(({row_reg, col_reg}==14'b00111011000000)) color_data = 12'b001000000100;
		if(({row_reg, col_reg}==14'b00111011000001)) color_data = 12'b001100000011;
		if(({row_reg, col_reg}==14'b00111011000010)) color_data = 12'b011100100011;
		if(({row_reg, col_reg}==14'b00111011000011)) color_data = 12'b100000110011;
		if(({row_reg, col_reg}==14'b00111011000100)) color_data = 12'b100001000011;
		if(({row_reg, col_reg}==14'b00111011000101)) color_data = 12'b101001100111;
		if(({row_reg, col_reg}==14'b00111011000110)) color_data = 12'b100101100111;
		if(({row_reg, col_reg}==14'b00111011000111)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}==14'b00111011001000)) color_data = 12'b001100010001;
		if(({row_reg, col_reg}>=14'b00111011001001) && ({row_reg, col_reg}<14'b00111011001011)) color_data = 12'b001100010010;
		if(({row_reg, col_reg}==14'b00111011001011)) color_data = 12'b001100010011;
		if(({row_reg, col_reg}>=14'b00111011001100) && ({row_reg, col_reg}<14'b00111011001110)) color_data = 12'b001100010010;
		if(({row_reg, col_reg}>=14'b00111011001110) && ({row_reg, col_reg}<14'b00111011010001)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}==14'b00111011010001)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}>=14'b00111011010010) && ({row_reg, col_reg}<14'b00111011010101)) color_data = 12'b010000100011;
		if(({row_reg, col_reg}>=14'b00111011010101) && ({row_reg, col_reg}<14'b00111011011000)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}==14'b00111011011000)) color_data = 12'b010000100011;
		if(({row_reg, col_reg}==14'b00111011011001)) color_data = 12'b001100010100;
		if(({row_reg, col_reg}==14'b00111011011010)) color_data = 12'b001000000101;
		if(({row_reg, col_reg}==14'b00111011011011)) color_data = 12'b000100000111;
		if(({row_reg, col_reg}==14'b00111011011100)) color_data = 12'b000000001010;
		if(({row_reg, col_reg}==14'b00111011011101)) color_data = 12'b000000001100;
		if(({row_reg, col_reg}==14'b00111011011110)) color_data = 12'b000000001110;

		if(({row_reg, col_reg}>=14'b00111011011111) && ({row_reg, col_reg}<14'b00111100111100)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=14'b00111100111100) && ({row_reg, col_reg}<14'b00111100111110)) color_data = 12'b000000001110;
		if(({row_reg, col_reg}==14'b00111100111110)) color_data = 12'b000000001101;
		if(({row_reg, col_reg}==14'b00111100111111)) color_data = 12'b000100001100;
		if(({row_reg, col_reg}==14'b00111101000000)) color_data = 12'b001000000100;
		if(({row_reg, col_reg}==14'b00111101000001)) color_data = 12'b001100000011;
		if(({row_reg, col_reg}==14'b00111101000010)) color_data = 12'b100001000110;
		if(({row_reg, col_reg}==14'b00111101000011)) color_data = 12'b110010001000;
		if(({row_reg, col_reg}==14'b00111101000100)) color_data = 12'b101110001000;
		if(({row_reg, col_reg}==14'b00111101000101)) color_data = 12'b101001110111;
		if(({row_reg, col_reg}==14'b00111101000110)) color_data = 12'b100101111000;
		if(({row_reg, col_reg}==14'b00111101000111)) color_data = 12'b011101010110;
		if(({row_reg, col_reg}==14'b00111101001000)) color_data = 12'b011101100111;
		if(({row_reg, col_reg}==14'b00111101001001)) color_data = 12'b010100110100;
		if(({row_reg, col_reg}==14'b00111101001010)) color_data = 12'b010000100011;
		if(({row_reg, col_reg}==14'b00111101001011)) color_data = 12'b010000100100;
		if(({row_reg, col_reg}>=14'b00111101001100) && ({row_reg, col_reg}<14'b00111101001110)) color_data = 12'b001100010011;
		if(({row_reg, col_reg}>=14'b00111101001110) && ({row_reg, col_reg}<14'b00111101010000)) color_data = 12'b001100100011;
		if(({row_reg, col_reg}==14'b00111101010000)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}==14'b00111101010001)) color_data = 12'b001100010010;
		if(({row_reg, col_reg}==14'b00111101010010)) color_data = 12'b001100100011;
		if(({row_reg, col_reg}>=14'b00111101010011) && ({row_reg, col_reg}<14'b00111101010111)) color_data = 12'b010000100011;
		if(({row_reg, col_reg}==14'b00111101010111)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}>=14'b00111101011000) && ({row_reg, col_reg}<14'b00111101011010)) color_data = 12'b010000100011;
		if(({row_reg, col_reg}==14'b00111101011010)) color_data = 12'b001100010100;
		if(({row_reg, col_reg}==14'b00111101011011)) color_data = 12'b001000010101;
		if(({row_reg, col_reg}==14'b00111101011100)) color_data = 12'b000100000111;
		if(({row_reg, col_reg}==14'b00111101011101)) color_data = 12'b000000001010;
		if(({row_reg, col_reg}==14'b00111101011110)) color_data = 12'b000000001101;

		if(({row_reg, col_reg}>=14'b00111101011111) && ({row_reg, col_reg}<14'b00111110111001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=14'b00111110111001) && ({row_reg, col_reg}<14'b00111110111101)) color_data = 12'b000000001110;
		if(({row_reg, col_reg}>=14'b00111110111101) && ({row_reg, col_reg}<14'b00111110111111)) color_data = 12'b000100001101;
		if(({row_reg, col_reg}==14'b00111110111111)) color_data = 12'b000100001100;
		if(({row_reg, col_reg}==14'b00111111000000)) color_data = 12'b000100000101;
		if(({row_reg, col_reg}==14'b00111111000001)) color_data = 12'b001000000100;
		if(({row_reg, col_reg}==14'b00111111000010)) color_data = 12'b100101101000;
		if(({row_reg, col_reg}==14'b00111111000011)) color_data = 12'b111110111100;
		if(({row_reg, col_reg}==14'b00111111000100)) color_data = 12'b110110101010;
		if(({row_reg, col_reg}>=14'b00111111000101) && ({row_reg, col_reg}<14'b00111111000111)) color_data = 12'b100101111000;
		if(({row_reg, col_reg}>=14'b00111111000111) && ({row_reg, col_reg}<14'b00111111001001)) color_data = 12'b100001111000;
		if(({row_reg, col_reg}==14'b00111111001001)) color_data = 12'b010000100100;
		if(({row_reg, col_reg}>=14'b00111111001010) && ({row_reg, col_reg}<14'b00111111001101)) color_data = 12'b000100000010;
		if(({row_reg, col_reg}==14'b00111111001101)) color_data = 12'b001000000010;
		if(({row_reg, col_reg}==14'b00111111001110)) color_data = 12'b001000010010;
		if(({row_reg, col_reg}==14'b00111111001111)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==14'b00111111010000)) color_data = 12'b001100010010;
		if(({row_reg, col_reg}>=14'b00111111010001) && ({row_reg, col_reg}<14'b00111111010110)) color_data = 12'b001100100011;
		if(({row_reg, col_reg}>=14'b00111111010110) && ({row_reg, col_reg}<14'b00111111011000)) color_data = 12'b010000100011;
		if(({row_reg, col_reg}>=14'b00111111011000) && ({row_reg, col_reg}<14'b00111111011010)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}==14'b00111111011010)) color_data = 12'b010000100011;
		if(({row_reg, col_reg}==14'b00111111011011)) color_data = 12'b001100010100;
		if(({row_reg, col_reg}==14'b00111111011100)) color_data = 12'b000100000101;
		if(({row_reg, col_reg}==14'b00111111011101)) color_data = 12'b000000001001;
		if(({row_reg, col_reg}==14'b00111111011110)) color_data = 12'b000000001100;

		if(({row_reg, col_reg}>=14'b00111111011111) && ({row_reg, col_reg}<14'b01000000110011)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==14'b01000000110011)) color_data = 12'b000000001110;
		if(({row_reg, col_reg}>=14'b01000000110100) && ({row_reg, col_reg}<14'b01000000111000)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==14'b01000000111000)) color_data = 12'b000100001110;
		if(({row_reg, col_reg}==14'b01000000111001)) color_data = 12'b001000001100;
		if(({row_reg, col_reg}==14'b01000000111010)) color_data = 12'b001100001010;
		if(({row_reg, col_reg}==14'b01000000111011)) color_data = 12'b010000001000;
		if(({row_reg, col_reg}==14'b01000000111100)) color_data = 12'b010100001000;
		if(({row_reg, col_reg}==14'b01000000111101)) color_data = 12'b010100000111;
		if(({row_reg, col_reg}==14'b01000000111110)) color_data = 12'b010000000111;
		if(({row_reg, col_reg}==14'b01000000111111)) color_data = 12'b010000001000;
		if(({row_reg, col_reg}==14'b01000001000000)) color_data = 12'b010000010011;
		if(({row_reg, col_reg}==14'b01000001000001)) color_data = 12'b010000000010;
		if(({row_reg, col_reg}==14'b01000001000010)) color_data = 12'b011001000100;
		if(({row_reg, col_reg}==14'b01000001000011)) color_data = 12'b100101110110;
		if(({row_reg, col_reg}==14'b01000001000100)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==14'b01000001000101)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==14'b01000001000110)) color_data = 12'b101010011010;
		if(({row_reg, col_reg}==14'b01000001000111)) color_data = 12'b100101111001;
		if(({row_reg, col_reg}==14'b01000001001000)) color_data = 12'b100001111010;
		if(({row_reg, col_reg}==14'b01000001001001)) color_data = 12'b010000111000;
		if(({row_reg, col_reg}==14'b01000001001010)) color_data = 12'b000100000111;
		if(({row_reg, col_reg}>=14'b01000001001011) && ({row_reg, col_reg}<14'b01000001001101)) color_data = 12'b000100001001;
		if(({row_reg, col_reg}==14'b01000001001101)) color_data = 12'b000100000110;
		if(({row_reg, col_reg}==14'b01000001001110)) color_data = 12'b000100000100;
		if(({row_reg, col_reg}==14'b01000001001111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==14'b01000001010000)) color_data = 12'b001100100011;
		if(({row_reg, col_reg}==14'b01000001010001)) color_data = 12'b001100010011;
		if(({row_reg, col_reg}==14'b01000001010010)) color_data = 12'b001100010010;
		if(({row_reg, col_reg}==14'b01000001010011)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}==14'b01000001010100)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==14'b01000001010101)) color_data = 12'b001100010010;
		if(({row_reg, col_reg}==14'b01000001010110)) color_data = 12'b010000010011;
		if(({row_reg, col_reg}==14'b01000001010111)) color_data = 12'b001100010100;
		if(({row_reg, col_reg}==14'b01000001011000)) color_data = 12'b010000010100;
		if(({row_reg, col_reg}==14'b01000001011001)) color_data = 12'b010000100011;
		if(({row_reg, col_reg}==14'b01000001011010)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==14'b01000001011011)) color_data = 12'b001100100011;
		if(({row_reg, col_reg}==14'b01000001011100)) color_data = 12'b001000010101;
		if(({row_reg, col_reg}==14'b01000001011101)) color_data = 12'b000000001000;
		if(({row_reg, col_reg}==14'b01000001011110)) color_data = 12'b000000001100;
		if(({row_reg, col_reg}==14'b01000001011111)) color_data = 12'b000000001110;

		if(({row_reg, col_reg}>=14'b01000001100000) && ({row_reg, col_reg}<14'b01000010110010)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==14'b01000010110010)) color_data = 12'b000000001110;
		if(({row_reg, col_reg}==14'b01000010110011)) color_data = 12'b000100001101;
		if(({row_reg, col_reg}>=14'b01000010110100) && ({row_reg, col_reg}<14'b01000010110110)) color_data = 12'b000100001110;
		if(({row_reg, col_reg}==14'b01000010110110)) color_data = 12'b000000001101;
		if(({row_reg, col_reg}==14'b01000010110111)) color_data = 12'b000100001101;
		if(({row_reg, col_reg}==14'b01000010111000)) color_data = 12'b001000001011;
		if(({row_reg, col_reg}==14'b01000010111001)) color_data = 12'b010000001001;
		if(({row_reg, col_reg}==14'b01000010111010)) color_data = 12'b010100001000;
		if(({row_reg, col_reg}==14'b01000010111011)) color_data = 12'b011100000111;
		if(({row_reg, col_reg}==14'b01000010111100)) color_data = 12'b100000010111;
		if(({row_reg, col_reg}==14'b01000010111101)) color_data = 12'b011100010110;
		if(({row_reg, col_reg}==14'b01000010111110)) color_data = 12'b011000000101;
		if(({row_reg, col_reg}==14'b01000010111111)) color_data = 12'b010100000101;
		if(({row_reg, col_reg}==14'b01000011000000)) color_data = 12'b010000000011;
		if(({row_reg, col_reg}==14'b01000011000001)) color_data = 12'b010000010010;
		if(({row_reg, col_reg}==14'b01000011000010)) color_data = 12'b010000010001;
		if(({row_reg, col_reg}==14'b01000011000011)) color_data = 12'b001100000001;
		if(({row_reg, col_reg}==14'b01000011000100)) color_data = 12'b011000110100;
		if(({row_reg, col_reg}==14'b01000011000101)) color_data = 12'b110010101011;
		if(({row_reg, col_reg}==14'b01000011000110)) color_data = 12'b110010101100;
		if(({row_reg, col_reg}==14'b01000011000111)) color_data = 12'b101010001010;
		if(({row_reg, col_reg}==14'b01000011001000)) color_data = 12'b100001011001;
		if(({row_reg, col_reg}==14'b01000011001001)) color_data = 12'b010100111000;
		if(({row_reg, col_reg}==14'b01000011001010)) color_data = 12'b001100011000;
		if(({row_reg, col_reg}>=14'b01000011001011) && ({row_reg, col_reg}<14'b01000011001101)) color_data = 12'b001000001001;
		if(({row_reg, col_reg}==14'b01000011001101)) color_data = 12'b000100000111;
		if(({row_reg, col_reg}==14'b01000011001110)) color_data = 12'b000100000101;
		if(({row_reg, col_reg}==14'b01000011001111)) color_data = 12'b000100000100;
		if(({row_reg, col_reg}==14'b01000011010000)) color_data = 12'b001000010101;
		if(({row_reg, col_reg}==14'b01000011010001)) color_data = 12'b001000010100;
		if(({row_reg, col_reg}==14'b01000011010010)) color_data = 12'b001100010011;
		if(({row_reg, col_reg}==14'b01000011010011)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}>=14'b01000011010100) && ({row_reg, col_reg}<14'b01000011010110)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}==14'b01000011010110)) color_data = 12'b001100010010;
		if(({row_reg, col_reg}>=14'b01000011010111) && ({row_reg, col_reg}<14'b01000011011001)) color_data = 12'b001100010011;
		if(({row_reg, col_reg}==14'b01000011011001)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==14'b01000011011010)) color_data = 12'b001100010010;
		if(({row_reg, col_reg}==14'b01000011011011)) color_data = 12'b001000010011;
		if(({row_reg, col_reg}==14'b01000011011100)) color_data = 12'b000100000101;
		if(({row_reg, col_reg}==14'b01000011011101)) color_data = 12'b000000001000;
		if(({row_reg, col_reg}==14'b01000011011110)) color_data = 12'b000000001100;

		if(({row_reg, col_reg}>=14'b01000011011111) && ({row_reg, col_reg}<14'b01000100110001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==14'b01000100110001)) color_data = 12'b000000001110;
		if(({row_reg, col_reg}==14'b01000100110010)) color_data = 12'b000100001101;
		if(({row_reg, col_reg}==14'b01000100110011)) color_data = 12'b001000001011;
		if(({row_reg, col_reg}>=14'b01000100110100) && ({row_reg, col_reg}<14'b01000100110110)) color_data = 12'b001100001010;
		if(({row_reg, col_reg}==14'b01000100110110)) color_data = 12'b001100001001;
		if(({row_reg, col_reg}==14'b01000100110111)) color_data = 12'b010000001001;
		if(({row_reg, col_reg}==14'b01000100111000)) color_data = 12'b011000001000;
		if(({row_reg, col_reg}==14'b01000100111001)) color_data = 12'b100000010111;
		if(({row_reg, col_reg}==14'b01000100111010)) color_data = 12'b101000100110;
		if(({row_reg, col_reg}>=14'b01000100111011) && ({row_reg, col_reg}<14'b01000100111101)) color_data = 12'b101100100110;
		if(({row_reg, col_reg}==14'b01000100111101)) color_data = 12'b101000100101;
		if(({row_reg, col_reg}>=14'b01000100111110) && ({row_reg, col_reg}<14'b01000101000000)) color_data = 12'b100000010100;
		if(({row_reg, col_reg}==14'b01000101000000)) color_data = 12'b011000000011;
		if(({row_reg, col_reg}==14'b01000101000001)) color_data = 12'b011000010011;
		if(({row_reg, col_reg}==14'b01000101000010)) color_data = 12'b010100010010;
		if(({row_reg, col_reg}==14'b01000101000011)) color_data = 12'b010000010010;
		if(({row_reg, col_reg}==14'b01000101000100)) color_data = 12'b011000110100;
		if(({row_reg, col_reg}==14'b01000101000101)) color_data = 12'b101110001001;
		if(({row_reg, col_reg}==14'b01000101000110)) color_data = 12'b101110001010;
		if(({row_reg, col_reg}==14'b01000101000111)) color_data = 12'b101001101001;
		if(({row_reg, col_reg}==14'b01000101001000)) color_data = 12'b100101011000;
		if(({row_reg, col_reg}==14'b01000101001001)) color_data = 12'b100001001000;
		if(({row_reg, col_reg}==14'b01000101001010)) color_data = 12'b011100101001;
		if(({row_reg, col_reg}==14'b01000101001011)) color_data = 12'b011000101001;
		if(({row_reg, col_reg}==14'b01000101001100)) color_data = 12'b010100011010;
		if(({row_reg, col_reg}==14'b01000101001101)) color_data = 12'b001100001001;
		if(({row_reg, col_reg}>=14'b01000101001110) && ({row_reg, col_reg}<14'b01000101010000)) color_data = 12'b000100001000;
		if(({row_reg, col_reg}==14'b01000101010000)) color_data = 12'b000000000111;
		if(({row_reg, col_reg}==14'b01000101010001)) color_data = 12'b000100000110;
		if(({row_reg, col_reg}==14'b01000101010010)) color_data = 12'b000100000101;
		if(({row_reg, col_reg}==14'b01000101010011)) color_data = 12'b001000000011;
		if(({row_reg, col_reg}==14'b01000101010100)) color_data = 12'b001100010011;
		if(({row_reg, col_reg}>=14'b01000101010101) && ({row_reg, col_reg}<14'b01000101010111)) color_data = 12'b001100010010;
		if(({row_reg, col_reg}>=14'b01000101010111) && ({row_reg, col_reg}<14'b01000101011001)) color_data = 12'b001100010011;
		if(({row_reg, col_reg}==14'b01000101011001)) color_data = 12'b001100100011;
		if(({row_reg, col_reg}==14'b01000101011010)) color_data = 12'b001100010100;
		if(({row_reg, col_reg}==14'b01000101011011)) color_data = 12'b001000000100;
		if(({row_reg, col_reg}==14'b01000101011100)) color_data = 12'b000100000111;
		if(({row_reg, col_reg}==14'b01000101011101)) color_data = 12'b000000001010;
		if(({row_reg, col_reg}==14'b01000101011110)) color_data = 12'b000000001110;

		if(({row_reg, col_reg}>=14'b01000101011111) && ({row_reg, col_reg}<14'b01000110101110)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=14'b01000110101110) && ({row_reg, col_reg}<14'b01000110110000)) color_data = 12'b000000001110;
		if(({row_reg, col_reg}==14'b01000110110000)) color_data = 12'b000000001101;
		if(({row_reg, col_reg}==14'b01000110110001)) color_data = 12'b000100001100;
		if(({row_reg, col_reg}==14'b01000110110010)) color_data = 12'b001100001010;
		if(({row_reg, col_reg}==14'b01000110110011)) color_data = 12'b010000001000;
		if(({row_reg, col_reg}==14'b01000110110100)) color_data = 12'b010100000111;
		if(({row_reg, col_reg}==14'b01000110110101)) color_data = 12'b011000010111;
		if(({row_reg, col_reg}==14'b01000110110110)) color_data = 12'b011100010110;
		if(({row_reg, col_reg}==14'b01000110110111)) color_data = 12'b100000010110;
		if(({row_reg, col_reg}==14'b01000110111000)) color_data = 12'b100100010101;
		if(({row_reg, col_reg}==14'b01000110111001)) color_data = 12'b101000100101;
		if(({row_reg, col_reg}>=14'b01000110111010) && ({row_reg, col_reg}<14'b01000110111101)) color_data = 12'b110000100100;
		if(({row_reg, col_reg}==14'b01000110111101)) color_data = 12'b101100010011;
		if(({row_reg, col_reg}>=14'b01000110111110) && ({row_reg, col_reg}<14'b01000111000000)) color_data = 12'b100100000010;
		if(({row_reg, col_reg}==14'b01000111000000)) color_data = 12'b100000010011;
		if(({row_reg, col_reg}==14'b01000111000001)) color_data = 12'b011000000010;
		if(({row_reg, col_reg}==14'b01000111000010)) color_data = 12'b011100010011;
		if(({row_reg, col_reg}==14'b01000111000011)) color_data = 12'b011100100100;
		if(({row_reg, col_reg}>=14'b01000111000100) && ({row_reg, col_reg}<14'b01000111000111)) color_data = 12'b010100010011;
		if(({row_reg, col_reg}==14'b01000111000111)) color_data = 12'b011000010100;
		if(({row_reg, col_reg}==14'b01000111001000)) color_data = 12'b011100010100;
		if(({row_reg, col_reg}==14'b01000111001001)) color_data = 12'b011100000100;
		if(({row_reg, col_reg}==14'b01000111001010)) color_data = 12'b011100000101;
		if(({row_reg, col_reg}==14'b01000111001011)) color_data = 12'b011100000110;
		if(({row_reg, col_reg}==14'b01000111001100)) color_data = 12'b011100011000;
		if(({row_reg, col_reg}==14'b01000111001101)) color_data = 12'b010100001000;
		if(({row_reg, col_reg}==14'b01000111001110)) color_data = 12'b001000001001;
		if(({row_reg, col_reg}==14'b01000111001111)) color_data = 12'b001000001010;
		if(({row_reg, col_reg}>=14'b01000111010000) && ({row_reg, col_reg}<14'b01000111010010)) color_data = 12'b000000001010;
		if(({row_reg, col_reg}==14'b01000111010010)) color_data = 12'b000100001000;
		if(({row_reg, col_reg}==14'b01000111010011)) color_data = 12'b000100000110;
		if(({row_reg, col_reg}==14'b01000111010100)) color_data = 12'b001000010101;
		if(({row_reg, col_reg}==14'b01000111010101)) color_data = 12'b001100010100;
		if(({row_reg, col_reg}==14'b01000111010110)) color_data = 12'b001100010011;
		if(({row_reg, col_reg}==14'b01000111010111)) color_data = 12'b001100010100;
		if(({row_reg, col_reg}==14'b01000111011000)) color_data = 12'b001000010100;
		if(({row_reg, col_reg}==14'b01000111011001)) color_data = 12'b001000010101;
		if(({row_reg, col_reg}==14'b01000111011010)) color_data = 12'b000100000101;
		if(({row_reg, col_reg}==14'b01000111011011)) color_data = 12'b000100000111;
		if(({row_reg, col_reg}==14'b01000111011100)) color_data = 12'b000000001010;
		if(({row_reg, col_reg}==14'b01000111011101)) color_data = 12'b000000001101;

		if(({row_reg, col_reg}>=14'b01000111011110) && ({row_reg, col_reg}<14'b01001000101101)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==14'b01001000101101)) color_data = 12'b000100001110;
		if(({row_reg, col_reg}==14'b01001000101110)) color_data = 12'b000100001100;
		if(({row_reg, col_reg}==14'b01001000101111)) color_data = 12'b001000001100;
		if(({row_reg, col_reg}==14'b01001000110000)) color_data = 12'b001100001010;
		if(({row_reg, col_reg}==14'b01001000110001)) color_data = 12'b010000001001;
		if(({row_reg, col_reg}==14'b01001000110010)) color_data = 12'b011000011000;
		if(({row_reg, col_reg}==14'b01001000110011)) color_data = 12'b100000100111;
		if(({row_reg, col_reg}==14'b01001000110100)) color_data = 12'b100100100110;
		if(({row_reg, col_reg}==14'b01001000110101)) color_data = 12'b101000100110;
		if(({row_reg, col_reg}==14'b01001000110110)) color_data = 12'b101000100101;
		if(({row_reg, col_reg}==14'b01001000110111)) color_data = 12'b101100100101;
		if(({row_reg, col_reg}==14'b01001000111000)) color_data = 12'b101100100100;
		if(({row_reg, col_reg}==14'b01001000111001)) color_data = 12'b110000100100;
		if(({row_reg, col_reg}>=14'b01001000111010) && ({row_reg, col_reg}<14'b01001000111100)) color_data = 12'b110000100011;
		if(({row_reg, col_reg}==14'b01001000111100)) color_data = 12'b110000100100;
		if(({row_reg, col_reg}==14'b01001000111101)) color_data = 12'b101100100011;
		if(({row_reg, col_reg}==14'b01001000111110)) color_data = 12'b100100010010;
		if(({row_reg, col_reg}==14'b01001000111111)) color_data = 12'b100100000010;
		if(({row_reg, col_reg}==14'b01001001000000)) color_data = 12'b100000010011;
		if(({row_reg, col_reg}>=14'b01001001000001) && ({row_reg, col_reg}<14'b01001001000011)) color_data = 12'b100000000011;
		if(({row_reg, col_reg}==14'b01001001000011)) color_data = 12'b100000010100;
		if(({row_reg, col_reg}==14'b01001001000100)) color_data = 12'b011000000011;
		if(({row_reg, col_reg}>=14'b01001001000101) && ({row_reg, col_reg}<14'b01001001000111)) color_data = 12'b010100000010;
		if(({row_reg, col_reg}==14'b01001001000111)) color_data = 12'b011100010011;
		if(({row_reg, col_reg}==14'b01001001001000)) color_data = 12'b100000010011;
		if(({row_reg, col_reg}>=14'b01001001001001) && ({row_reg, col_reg}<14'b01001001001011)) color_data = 12'b100100000011;
		if(({row_reg, col_reg}==14'b01001001001011)) color_data = 12'b100100010011;
		if(({row_reg, col_reg}==14'b01001001001100)) color_data = 12'b100100100101;
		if(({row_reg, col_reg}==14'b01001001001101)) color_data = 12'b011100010111;
		if(({row_reg, col_reg}==14'b01001001001110)) color_data = 12'b010000001000;
		if(({row_reg, col_reg}==14'b01001001001111)) color_data = 12'b001100001001;
		if(({row_reg, col_reg}>=14'b01001001010000) && ({row_reg, col_reg}<14'b01001001010010)) color_data = 12'b000000001100;
		if(({row_reg, col_reg}==14'b01001001010010)) color_data = 12'b000000001011;
		if(({row_reg, col_reg}==14'b01001001010011)) color_data = 12'b000000001001;
		if(({row_reg, col_reg}==14'b01001001010100)) color_data = 12'b000000001000;
		if(({row_reg, col_reg}==14'b01001001010101)) color_data = 12'b000000000110;
		if(({row_reg, col_reg}>=14'b01001001010110) && ({row_reg, col_reg}<14'b01001001011000)) color_data = 12'b000000000101;
		if(({row_reg, col_reg}==14'b01001001011000)) color_data = 12'b000100000110;
		if(({row_reg, col_reg}==14'b01001001011001)) color_data = 12'b000000000111;
		if(({row_reg, col_reg}==14'b01001001011010)) color_data = 12'b000000001000;
		if(({row_reg, col_reg}==14'b01001001011011)) color_data = 12'b000000001010;
		if(({row_reg, col_reg}==14'b01001001011100)) color_data = 12'b000000001101;
		if(({row_reg, col_reg}==14'b01001001011101)) color_data = 12'b000000001110;

		if(({row_reg, col_reg}>=14'b01001001011110) && ({row_reg, col_reg}<14'b01001010101100)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==14'b01001010101100)) color_data = 12'b000100001101;
		if(({row_reg, col_reg}==14'b01001010101101)) color_data = 12'b001000001100;
		if(({row_reg, col_reg}==14'b01001010101110)) color_data = 12'b001100001010;
		if(({row_reg, col_reg}==14'b01001010101111)) color_data = 12'b010000001010;
		if(({row_reg, col_reg}==14'b01001010110000)) color_data = 12'b011000000111;
		if(({row_reg, col_reg}==14'b01001010110001)) color_data = 12'b011100010111;
		if(({row_reg, col_reg}==14'b01001010110010)) color_data = 12'b100100010110;
		if(({row_reg, col_reg}==14'b01001010110011)) color_data = 12'b101000100101;
		if(({row_reg, col_reg}==14'b01001010110100)) color_data = 12'b101100100100;
		if(({row_reg, col_reg}>=14'b01001010110101) && ({row_reg, col_reg}<14'b01001010110111)) color_data = 12'b101000010010;
		if(({row_reg, col_reg}==14'b01001010110111)) color_data = 12'b101100100100;
		if(({row_reg, col_reg}>=14'b01001010111000) && ({row_reg, col_reg}<14'b01001010111011)) color_data = 12'b110000100100;
		if(({row_reg, col_reg}==14'b01001010111011)) color_data = 12'b101100010011;
		if(({row_reg, col_reg}==14'b01001010111100)) color_data = 12'b101000000011;
		if(({row_reg, col_reg}==14'b01001010111101)) color_data = 12'b101000010011;
		if(({row_reg, col_reg}==14'b01001010111110)) color_data = 12'b101000010100;
		if(({row_reg, col_reg}==14'b01001010111111)) color_data = 12'b101000100100;
		if(({row_reg, col_reg}==14'b01001011000000)) color_data = 12'b101000010011;
		if(({row_reg, col_reg}==14'b01001011000001)) color_data = 12'b101100100101;
		if(({row_reg, col_reg}==14'b01001011000010)) color_data = 12'b100100010100;
		if(({row_reg, col_reg}>=14'b01001011000011) && ({row_reg, col_reg}<14'b01001011000101)) color_data = 12'b100000000100;
		if(({row_reg, col_reg}==14'b01001011000101)) color_data = 12'b100000010100;
		if(({row_reg, col_reg}==14'b01001011000110)) color_data = 12'b011100000011;
		if(({row_reg, col_reg}==14'b01001011000111)) color_data = 12'b100100100100;
		if(({row_reg, col_reg}==14'b01001011001000)) color_data = 12'b101000100100;
		if(({row_reg, col_reg}==14'b01001011001001)) color_data = 12'b101100100100;
		if(({row_reg, col_reg}==14'b01001011001010)) color_data = 12'b101100010011;
		if(({row_reg, col_reg}==14'b01001011001011)) color_data = 12'b101100100011;
		if(({row_reg, col_reg}==14'b01001011001100)) color_data = 12'b101100100100;
		if(({row_reg, col_reg}==14'b01001011001101)) color_data = 12'b101000110110;
		if(({row_reg, col_reg}==14'b01001011001110)) color_data = 12'b100000100111;
		if(({row_reg, col_reg}==14'b01001011001111)) color_data = 12'b010100000110;
		if(({row_reg, col_reg}>=14'b01001011010000) && ({row_reg, col_reg}<14'b01001011010010)) color_data = 12'b000100001101;
		if(({row_reg, col_reg}>=14'b01001011010010) && ({row_reg, col_reg}<14'b01001011010100)) color_data = 12'b000000001101;
		if(({row_reg, col_reg}==14'b01001011010100)) color_data = 12'b000000001100;
		if(({row_reg, col_reg}==14'b01001011010101)) color_data = 12'b000000001011;
		if(({row_reg, col_reg}>=14'b01001011010110) && ({row_reg, col_reg}<14'b01001011011001)) color_data = 12'b000000001010;
		if(({row_reg, col_reg}==14'b01001011011001)) color_data = 12'b000000001011;
		if(({row_reg, col_reg}==14'b01001011011010)) color_data = 12'b000000001100;
		if(({row_reg, col_reg}==14'b01001011011011)) color_data = 12'b000000001101;

		if(({row_reg, col_reg}>=14'b01001011011100) && ({row_reg, col_reg}<14'b01001100101011)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==14'b01001100101011)) color_data = 12'b000000001101;
		if(({row_reg, col_reg}==14'b01001100101100)) color_data = 12'b001000001100;
		if(({row_reg, col_reg}==14'b01001100101101)) color_data = 12'b010000001001;
		if(({row_reg, col_reg}==14'b01001100101110)) color_data = 12'b010100001000;
		if(({row_reg, col_reg}==14'b01001100101111)) color_data = 12'b011000011000;
		if(({row_reg, col_reg}==14'b01001100110000)) color_data = 12'b100100100110;
		if(({row_reg, col_reg}==14'b01001100110001)) color_data = 12'b101000100110;
		if(({row_reg, col_reg}==14'b01001100110010)) color_data = 12'b101100110101;
		if(({row_reg, col_reg}==14'b01001100110011)) color_data = 12'b110000100100;
		if(({row_reg, col_reg}==14'b01001100110100)) color_data = 12'b101100010011;
		if(({row_reg, col_reg}==14'b01001100110101)) color_data = 12'b100100000001;
		if(({row_reg, col_reg}==14'b01001100110110)) color_data = 12'b101000000010;
		if(({row_reg, col_reg}>=14'b01001100110111) && ({row_reg, col_reg}<14'b01001100111010)) color_data = 12'b110000100100;
		if(({row_reg, col_reg}==14'b01001100111010)) color_data = 12'b110000100101;
		if(({row_reg, col_reg}==14'b01001100111011)) color_data = 12'b101100010100;
		if(({row_reg, col_reg}>=14'b01001100111100) && ({row_reg, col_reg}<14'b01001100111110)) color_data = 12'b100100000011;
		if(({row_reg, col_reg}==14'b01001100111110)) color_data = 12'b101100100101;
		if(({row_reg, col_reg}==14'b01001100111111)) color_data = 12'b101100110110;
		if(({row_reg, col_reg}==14'b01001101000000)) color_data = 12'b101100100100;
		if(({row_reg, col_reg}==14'b01001101000001)) color_data = 12'b110000110110;
		if(({row_reg, col_reg}==14'b01001101000010)) color_data = 12'b101000010100;
		if(({row_reg, col_reg}==14'b01001101000011)) color_data = 12'b100100000100;
		if(({row_reg, col_reg}>=14'b01001101000100) && ({row_reg, col_reg}<14'b01001101000110)) color_data = 12'b100000000100;
		if(({row_reg, col_reg}==14'b01001101000110)) color_data = 12'b100000000011;
		if(({row_reg, col_reg}==14'b01001101000111)) color_data = 12'b101000110101;
		if(({row_reg, col_reg}==14'b01001101001000)) color_data = 12'b101100110101;
		if(({row_reg, col_reg}==14'b01001101001001)) color_data = 12'b110000110101;
		if(({row_reg, col_reg}==14'b01001101001010)) color_data = 12'b110000100100;
		if(({row_reg, col_reg}>=14'b01001101001011) && ({row_reg, col_reg}<14'b01001101001101)) color_data = 12'b110000100011;
		if(({row_reg, col_reg}==14'b01001101001101)) color_data = 12'b101100100100;
		if(({row_reg, col_reg}==14'b01001101001110)) color_data = 12'b101000100101;
		if(({row_reg, col_reg}==14'b01001101001111)) color_data = 12'b011100000100;
		if(({row_reg, col_reg}==14'b01001101010000)) color_data = 12'b010000001011;
		if(({row_reg, col_reg}==14'b01001101010001)) color_data = 12'b001000001011;
		if(({row_reg, col_reg}==14'b01001101010010)) color_data = 12'b000100001101;
		if(({row_reg, col_reg}>=14'b01001101010011) && ({row_reg, col_reg}<14'b01001101011000)) color_data = 12'b000000001110;
		if(({row_reg, col_reg}==14'b01001101011000)) color_data = 12'b000000001101;
		if(({row_reg, col_reg}>=14'b01001101011001) && ({row_reg, col_reg}<14'b01001101011011)) color_data = 12'b000000001110;

		if(({row_reg, col_reg}>=14'b01001101011011) && ({row_reg, col_reg}<14'b01001110101010)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==14'b01001110101010)) color_data = 12'b000000001110;
		if(({row_reg, col_reg}==14'b01001110101011)) color_data = 12'b000100001100;
		if(({row_reg, col_reg}==14'b01001110101100)) color_data = 12'b001100001010;
		if(({row_reg, col_reg}==14'b01001110101101)) color_data = 12'b010100000111;
		if(({row_reg, col_reg}==14'b01001110101110)) color_data = 12'b011100010110;
		if(({row_reg, col_reg}==14'b01001110101111)) color_data = 12'b100100100101;
		if(({row_reg, col_reg}==14'b01001110110000)) color_data = 12'b100100010100;
		if(({row_reg, col_reg}==14'b01001110110001)) color_data = 12'b100100010011;
		if(({row_reg, col_reg}>=14'b01001110110010) && ({row_reg, col_reg}<14'b01001110110101)) color_data = 12'b101000010011;
		if(({row_reg, col_reg}==14'b01001110110101)) color_data = 12'b100100000010;
		if(({row_reg, col_reg}==14'b01001110110110)) color_data = 12'b100100000011;
		if(({row_reg, col_reg}==14'b01001110110111)) color_data = 12'b101000010011;
		if(({row_reg, col_reg}==14'b01001110111000)) color_data = 12'b101000010100;
		if(({row_reg, col_reg}==14'b01001110111001)) color_data = 12'b100100010011;
		if(({row_reg, col_reg}==14'b01001110111010)) color_data = 12'b101000010100;
		if(({row_reg, col_reg}==14'b01001110111011)) color_data = 12'b101000010011;
		if(({row_reg, col_reg}==14'b01001110111100)) color_data = 12'b100000000010;
		if(({row_reg, col_reg}==14'b01001110111101)) color_data = 12'b100100000011;
		if(({row_reg, col_reg}>=14'b01001110111110) && ({row_reg, col_reg}<14'b01001111000000)) color_data = 12'b101000010100;
		if(({row_reg, col_reg}==14'b01001111000000)) color_data = 12'b101000010011;
		if(({row_reg, col_reg}==14'b01001111000001)) color_data = 12'b101000010100;
		if(({row_reg, col_reg}>=14'b01001111000010) && ({row_reg, col_reg}<14'b01001111000101)) color_data = 12'b100100000100;
		if(({row_reg, col_reg}>=14'b01001111000101) && ({row_reg, col_reg}<14'b01001111000111)) color_data = 12'b100000000011;
		if(({row_reg, col_reg}==14'b01001111000111)) color_data = 12'b100100010100;
		if(({row_reg, col_reg}>=14'b01001111001000) && ({row_reg, col_reg}<14'b01001111001010)) color_data = 12'b101000010100;
		if(({row_reg, col_reg}==14'b01001111001010)) color_data = 12'b101100010011;
		if(({row_reg, col_reg}==14'b01001111001011)) color_data = 12'b110000010100;
		if(({row_reg, col_reg}==14'b01001111001100)) color_data = 12'b110000010011;
		if(({row_reg, col_reg}==14'b01001111001101)) color_data = 12'b110000100100;
		if(({row_reg, col_reg}==14'b01001111001110)) color_data = 12'b110000100101;
		if(({row_reg, col_reg}==14'b01001111001111)) color_data = 12'b101100100101;
		if(({row_reg, col_reg}==14'b01001111010000)) color_data = 12'b100000101001;
		if(({row_reg, col_reg}==14'b01001111010001)) color_data = 12'b010100001001;
		if(({row_reg, col_reg}==14'b01001111010010)) color_data = 12'b001100001011;
		if(({row_reg, col_reg}==14'b01001111010011)) color_data = 12'b000100001101;
		if(({row_reg, col_reg}>=14'b01001111010100) && ({row_reg, col_reg}<14'b01001111011010)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==14'b01001111011010)) color_data = 12'b000000001110;

		if(({row_reg, col_reg}>=14'b01001111011011) && ({row_reg, col_reg}<14'b01010000101010)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==14'b01010000101010)) color_data = 12'b000100001101;
		if(({row_reg, col_reg}==14'b01010000101011)) color_data = 12'b001000001011;
		if(({row_reg, col_reg}==14'b01010000101100)) color_data = 12'b010000001000;
		if(({row_reg, col_reg}==14'b01010000101101)) color_data = 12'b100000010111;
		if(({row_reg, col_reg}==14'b01010000101110)) color_data = 12'b011100000011;
		if(({row_reg, col_reg}==14'b01010000101111)) color_data = 12'b100000000010;
		if(({row_reg, col_reg}==14'b01010000110000)) color_data = 12'b100000010011;
		if(({row_reg, col_reg}>=14'b01010000110001) && ({row_reg, col_reg}<14'b01010000110011)) color_data = 12'b100000000010;
		if(({row_reg, col_reg}>=14'b01010000110011) && ({row_reg, col_reg}<14'b01010000110110)) color_data = 12'b100000000011;
		if(({row_reg, col_reg}==14'b01010000110110)) color_data = 12'b100000010100;
		if(({row_reg, col_reg}==14'b01010000110111)) color_data = 12'b011100000011;
		if(({row_reg, col_reg}==14'b01010000111000)) color_data = 12'b100000000011;
		if(({row_reg, col_reg}==14'b01010000111001)) color_data = 12'b100000010011;
		if(({row_reg, col_reg}==14'b01010000111010)) color_data = 12'b100000000010;
		if(({row_reg, col_reg}>=14'b01010000111011) && ({row_reg, col_reg}<14'b01010000111111)) color_data = 12'b100000000011;
		if(({row_reg, col_reg}==14'b01010000111111)) color_data = 12'b100000000010;
		if(({row_reg, col_reg}==14'b01010001000000)) color_data = 12'b011100000010;
		if(({row_reg, col_reg}>=14'b01010001000001) && ({row_reg, col_reg}<14'b01010001000011)) color_data = 12'b100000000011;
		if(({row_reg, col_reg}>=14'b01010001000011) && ({row_reg, col_reg}<14'b01010001000101)) color_data = 12'b100100000100;
		if(({row_reg, col_reg}==14'b01010001000101)) color_data = 12'b100100000011;
		if(({row_reg, col_reg}==14'b01010001000110)) color_data = 12'b100000000011;
		if(({row_reg, col_reg}==14'b01010001000111)) color_data = 12'b100000000010;
		if(({row_reg, col_reg}>=14'b01010001001000) && ({row_reg, col_reg}<14'b01010001001010)) color_data = 12'b100000000011;
		if(({row_reg, col_reg}==14'b01010001001010)) color_data = 12'b100100000011;
		if(({row_reg, col_reg}==14'b01010001001011)) color_data = 12'b101000010100;
		if(({row_reg, col_reg}>=14'b01010001001100) && ({row_reg, col_reg}<14'b01010001001110)) color_data = 12'b110000100101;
		if(({row_reg, col_reg}>=14'b01010001001110) && ({row_reg, col_reg}<14'b01010001010000)) color_data = 12'b110000100100;
		if(({row_reg, col_reg}==14'b01010001010000)) color_data = 12'b101000100110;
		if(({row_reg, col_reg}==14'b01010001010001)) color_data = 12'b011100000110;
		if(({row_reg, col_reg}==14'b01010001010010)) color_data = 12'b010000001000;
		if(({row_reg, col_reg}==14'b01010001010011)) color_data = 12'b001000001011;
		if(({row_reg, col_reg}==14'b01010001010100)) color_data = 12'b000000001101;

		if(({row_reg, col_reg}>=14'b01010001010101) && ({row_reg, col_reg}<14'b01010010101010)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==14'b01010010101010)) color_data = 12'b000100001101;
		if(({row_reg, col_reg}==14'b01010010101011)) color_data = 12'b001100001010;
		if(({row_reg, col_reg}==14'b01010010101100)) color_data = 12'b010100000111;
		if(({row_reg, col_reg}==14'b01010010101101)) color_data = 12'b100000010110;
		if(({row_reg, col_reg}==14'b01010010101110)) color_data = 12'b100000000011;
		if(({row_reg, col_reg}==14'b01010010101111)) color_data = 12'b100100010010;
		if(({row_reg, col_reg}>=14'b01010010110000) && ({row_reg, col_reg}<14'b01010010110011)) color_data = 12'b011100010011;
		if(({row_reg, col_reg}>=14'b01010010110011) && ({row_reg, col_reg}<14'b01010010110101)) color_data = 12'b011100010100;
		if(({row_reg, col_reg}==14'b01010010110101)) color_data = 12'b011000010011;
		if(({row_reg, col_reg}==14'b01010010110110)) color_data = 12'b011000010100;
		if(({row_reg, col_reg}>=14'b01010010110111) && ({row_reg, col_reg}<14'b01010010111001)) color_data = 12'b011000010011;
		if(({row_reg, col_reg}==14'b01010010111001)) color_data = 12'b011100010011;
		if(({row_reg, col_reg}==14'b01010010111010)) color_data = 12'b011000010011;
		if(({row_reg, col_reg}==14'b01010010111011)) color_data = 12'b011100010011;
		if(({row_reg, col_reg}==14'b01010010111100)) color_data = 12'b100000100101;
		if(({row_reg, col_reg}>=14'b01010010111101) && ({row_reg, col_reg}<14'b01010011000001)) color_data = 12'b100000100100;
		if(({row_reg, col_reg}==14'b01010011000001)) color_data = 12'b100000100101;
		if(({row_reg, col_reg}==14'b01010011000010)) color_data = 12'b011100010011;
		if(({row_reg, col_reg}>=14'b01010011000011) && ({row_reg, col_reg}<14'b01010011000111)) color_data = 12'b100000000011;
		if(({row_reg, col_reg}==14'b01010011000111)) color_data = 12'b100100010100;
		if(({row_reg, col_reg}>=14'b01010011001000) && ({row_reg, col_reg}<14'b01010011001011)) color_data = 12'b100000000011;
		if(({row_reg, col_reg}==14'b01010011001011)) color_data = 12'b100100010100;
		if(({row_reg, col_reg}==14'b01010011001100)) color_data = 12'b101000010101;
		if(({row_reg, col_reg}==14'b01010011001101)) color_data = 12'b101100010101;
		if(({row_reg, col_reg}==14'b01010011001110)) color_data = 12'b101100010100;
		if(({row_reg, col_reg}==14'b01010011001111)) color_data = 12'b101100100100;
		if(({row_reg, col_reg}==14'b01010011010000)) color_data = 12'b101100100011;
		if(({row_reg, col_reg}==14'b01010011010001)) color_data = 12'b101000010101;
		if(({row_reg, col_reg}==14'b01010011010010)) color_data = 12'b011100010111;
		if(({row_reg, col_reg}==14'b01010011010011)) color_data = 12'b010000001001;
		if(({row_reg, col_reg}==14'b01010011010100)) color_data = 12'b001000001011;
		if(({row_reg, col_reg}==14'b01010011010101)) color_data = 12'b000100001101;
		if(({row_reg, col_reg}==14'b01010011010110)) color_data = 12'b000000001110;

		if(({row_reg, col_reg}>=14'b01010011010111) && ({row_reg, col_reg}<14'b01010100101001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==14'b01010100101001)) color_data = 12'b000000001110;
		if(({row_reg, col_reg}==14'b01010100101010)) color_data = 12'b000100001101;
		if(({row_reg, col_reg}==14'b01010100101011)) color_data = 12'b001100001010;
		if(({row_reg, col_reg}==14'b01010100101100)) color_data = 12'b010100000111;
		if(({row_reg, col_reg}==14'b01010100101101)) color_data = 12'b100000010101;
		if(({row_reg, col_reg}==14'b01010100101110)) color_data = 12'b100000000010;
		if(({row_reg, col_reg}==14'b01010100101111)) color_data = 12'b100000010010;
		if(({row_reg, col_reg}>=14'b01010100110000) && ({row_reg, col_reg}<14'b01010100110010)) color_data = 12'b011100100100;
		if(({row_reg, col_reg}==14'b01010100110010)) color_data = 12'b011100100101;
		if(({row_reg, col_reg}==14'b01010100110011)) color_data = 12'b011100110101;
		if(({row_reg, col_reg}==14'b01010100110100)) color_data = 12'b011000100100;
		if(({row_reg, col_reg}==14'b01010100110101)) color_data = 12'b010000010011;
		if(({row_reg, col_reg}==14'b01010100110110)) color_data = 12'b010000000010;
		if(({row_reg, col_reg}==14'b01010100110111)) color_data = 12'b010000010011;
		if(({row_reg, col_reg}==14'b01010100111000)) color_data = 12'b010100010011;
		if(({row_reg, col_reg}==14'b01010100111001)) color_data = 12'b010000010010;
		if(({row_reg, col_reg}==14'b01010100111010)) color_data = 12'b010000000010;
		if(({row_reg, col_reg}==14'b01010100111011)) color_data = 12'b011100110101;
		if(({row_reg, col_reg}==14'b01010100111100)) color_data = 12'b101001111001;
		if(({row_reg, col_reg}==14'b01010100111101)) color_data = 12'b101101111001;
		if(({row_reg, col_reg}==14'b01010100111110)) color_data = 12'b101001111001;
		if(({row_reg, col_reg}>=14'b01010100111111) && ({row_reg, col_reg}<14'b01010101000010)) color_data = 12'b101101111001;
		if(({row_reg, col_reg}==14'b01010101000010)) color_data = 12'b100101000101;
		if(({row_reg, col_reg}==14'b01010101000011)) color_data = 12'b011100100011;
		if(({row_reg, col_reg}==14'b01010101000100)) color_data = 12'b011100010011;
		if(({row_reg, col_reg}==14'b01010101000101)) color_data = 12'b100000010011;
		if(({row_reg, col_reg}>=14'b01010101000110) && ({row_reg, col_reg}<14'b01010101001000)) color_data = 12'b011100000011;
		if(({row_reg, col_reg}==14'b01010101001000)) color_data = 12'b100000010100;
		if(({row_reg, col_reg}==14'b01010101001001)) color_data = 12'b011100000011;
		if(({row_reg, col_reg}==14'b01010101001010)) color_data = 12'b011100010011;
		if(({row_reg, col_reg}==14'b01010101001011)) color_data = 12'b100000010011;
		if(({row_reg, col_reg}>=14'b01010101001100) && ({row_reg, col_reg}<14'b01010101001111)) color_data = 12'b100000000011;
		if(({row_reg, col_reg}==14'b01010101001111)) color_data = 12'b100000000010;
		if(({row_reg, col_reg}==14'b01010101010000)) color_data = 12'b101100100011;
		if(({row_reg, col_reg}==14'b01010101010001)) color_data = 12'b101100100100;
		if(({row_reg, col_reg}==14'b01010101010010)) color_data = 12'b101000100111;
		if(({row_reg, col_reg}==14'b01010101010011)) color_data = 12'b011100011000;
		if(({row_reg, col_reg}==14'b01010101010100)) color_data = 12'b010000001001;
		if(({row_reg, col_reg}==14'b01010101010101)) color_data = 12'b001000001011;
		if(({row_reg, col_reg}==14'b01010101010110)) color_data = 12'b000100001101;

		if(({row_reg, col_reg}>=14'b01010101010111) && ({row_reg, col_reg}<14'b01010110101001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==14'b01010110101001)) color_data = 12'b000000001110;
		if(({row_reg, col_reg}==14'b01010110101010)) color_data = 12'b000100001100;
		if(({row_reg, col_reg}==14'b01010110101011)) color_data = 12'b001100001001;
		if(({row_reg, col_reg}==14'b01010110101100)) color_data = 12'b010100000110;
		if(({row_reg, col_reg}==14'b01010110101101)) color_data = 12'b011100010101;
		if(({row_reg, col_reg}>=14'b01010110101110) && ({row_reg, col_reg}<14'b01010110110000)) color_data = 12'b011100010011;
		if(({row_reg, col_reg}>=14'b01010110110000) && ({row_reg, col_reg}<14'b01010110110100)) color_data = 12'b011000110100;
		if(({row_reg, col_reg}==14'b01010110110100)) color_data = 12'b010100100011;
		if(({row_reg, col_reg}==14'b01010110110101)) color_data = 12'b010000010010;
		if(({row_reg, col_reg}==14'b01010110110110)) color_data = 12'b001100010010;
		if(({row_reg, col_reg}==14'b01010110110111)) color_data = 12'b010000010011;
		if(({row_reg, col_reg}==14'b01010110111000)) color_data = 12'b001100010010;
		if(({row_reg, col_reg}==14'b01010110111001)) color_data = 12'b010000010010;
		if(({row_reg, col_reg}==14'b01010110111010)) color_data = 12'b010000010011;
		if(({row_reg, col_reg}==14'b01010110111011)) color_data = 12'b011001000101;
		if(({row_reg, col_reg}>=14'b01010110111100) && ({row_reg, col_reg}<14'b01010110111110)) color_data = 12'b101010001001;
		if(({row_reg, col_reg}>=14'b01010110111110) && ({row_reg, col_reg}<14'b01010111000000)) color_data = 12'b100101111000;
		if(({row_reg, col_reg}==14'b01010111000000)) color_data = 12'b101001111001;
		if(({row_reg, col_reg}==14'b01010111000001)) color_data = 12'b101110001001;
		if(({row_reg, col_reg}==14'b01010111000010)) color_data = 12'b100001000101;
		if(({row_reg, col_reg}==14'b01010111000011)) color_data = 12'b010100010010;
		if(({row_reg, col_reg}==14'b01010111000100)) color_data = 12'b011000010011;
		if(({row_reg, col_reg}==14'b01010111000101)) color_data = 12'b100000100101;
		if(({row_reg, col_reg}>=14'b01010111000110) && ({row_reg, col_reg}<14'b01010111001001)) color_data = 12'b011100010100;
		if(({row_reg, col_reg}>=14'b01010111001001) && ({row_reg, col_reg}<14'b01010111001101)) color_data = 12'b011100010011;
		if(({row_reg, col_reg}>=14'b01010111001101) && ({row_reg, col_reg}<14'b01010111010000)) color_data = 12'b100000010011;
		if(({row_reg, col_reg}==14'b01010111010000)) color_data = 12'b101100100011;
		if(({row_reg, col_reg}==14'b01010111010001)) color_data = 12'b101100100100;
		if(({row_reg, col_reg}==14'b01010111010010)) color_data = 12'b101100100101;
		if(({row_reg, col_reg}==14'b01010111010011)) color_data = 12'b100100100111;
		if(({row_reg, col_reg}==14'b01010111010100)) color_data = 12'b011100000111;
		if(({row_reg, col_reg}==14'b01010111010101)) color_data = 12'b010000001001;
		if(({row_reg, col_reg}==14'b01010111010110)) color_data = 12'b001000001011;
		if(({row_reg, col_reg}==14'b01010111010111)) color_data = 12'b000000001110;

		if(({row_reg, col_reg}>=14'b01010111011000) && ({row_reg, col_reg}<14'b01011000101001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==14'b01011000101001)) color_data = 12'b000000001101;
		if(({row_reg, col_reg}==14'b01011000101010)) color_data = 12'b000100001011;
		if(({row_reg, col_reg}==14'b01011000101011)) color_data = 12'b001100001000;
		if(({row_reg, col_reg}==14'b01011000101100)) color_data = 12'b010000000101;
		if(({row_reg, col_reg}==14'b01011000101101)) color_data = 12'b011100010101;
		if(({row_reg, col_reg}>=14'b01011000101110) && ({row_reg, col_reg}<14'b01011000110000)) color_data = 12'b011100100100;
		if(({row_reg, col_reg}==14'b01011000110000)) color_data = 12'b010100110100;
		if(({row_reg, col_reg}==14'b01011000110001)) color_data = 12'b010100110011;
		if(({row_reg, col_reg}>=14'b01011000110010) && ({row_reg, col_reg}<14'b01011000110100)) color_data = 12'b011000110100;
		if(({row_reg, col_reg}==14'b01011000110100)) color_data = 12'b010100100011;
		if(({row_reg, col_reg}==14'b01011000110101)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}==14'b01011000110110)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==14'b01011000110111)) color_data = 12'b001100010010;
		if(({row_reg, col_reg}==14'b01011000111000)) color_data = 12'b010000100011;
		if(({row_reg, col_reg}==14'b01011000111001)) color_data = 12'b011101010110;
		if(({row_reg, col_reg}==14'b01011000111010)) color_data = 12'b100001100111;
		if(({row_reg, col_reg}==14'b01011000111011)) color_data = 12'b100101111000;
		if(({row_reg, col_reg}==14'b01011000111100)) color_data = 12'b101010001001;
		if(({row_reg, col_reg}>=14'b01011000111101) && ({row_reg, col_reg}<14'b01011001000000)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==14'b01011001000000)) color_data = 12'b100101111000;
		if(({row_reg, col_reg}==14'b01011001000001)) color_data = 12'b101010001000;
		if(({row_reg, col_reg}==14'b01011001000010)) color_data = 12'b011101000100;
		if(({row_reg, col_reg}==14'b01011001000011)) color_data = 12'b001100000001;
		if(({row_reg, col_reg}==14'b01011001000100)) color_data = 12'b011000100011;
		if(({row_reg, col_reg}==14'b01011001000101)) color_data = 12'b101001101000;
		if(({row_reg, col_reg}==14'b01011001000110)) color_data = 12'b101001011000;
		if(({row_reg, col_reg}>=14'b01011001000111) && ({row_reg, col_reg}<14'b01011001001010)) color_data = 12'b101001101000;
		if(({row_reg, col_reg}>=14'b01011001001010) && ({row_reg, col_reg}<14'b01011001001100)) color_data = 12'b101001100111;
		if(({row_reg, col_reg}==14'b01011001001100)) color_data = 12'b101001010111;
		if(({row_reg, col_reg}>=14'b01011001001101) && ({row_reg, col_reg}<14'b01011001010000)) color_data = 12'b101001100111;
		if(({row_reg, col_reg}==14'b01011001010000)) color_data = 12'b101000100011;
		if(({row_reg, col_reg}==14'b01011001010001)) color_data = 12'b100100000010;
		if(({row_reg, col_reg}==14'b01011001010010)) color_data = 12'b101000010100;
		if(({row_reg, col_reg}==14'b01011001010011)) color_data = 12'b101100100110;
		if(({row_reg, col_reg}==14'b01011001010100)) color_data = 12'b100100100111;
		if(({row_reg, col_reg}==14'b01011001010101)) color_data = 12'b011000011000;
		if(({row_reg, col_reg}==14'b01011001010110)) color_data = 12'b001100001010;
		if(({row_reg, col_reg}==14'b01011001010111)) color_data = 12'b000100001100;

		if(({row_reg, col_reg}>=14'b01011001011000) && ({row_reg, col_reg}<14'b01011010101000)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==14'b01011010101000)) color_data = 12'b000000001110;
		if(({row_reg, col_reg}==14'b01011010101001)) color_data = 12'b000100001100;
		if(({row_reg, col_reg}==14'b01011010101010)) color_data = 12'b000100001001;
		if(({row_reg, col_reg}==14'b01011010101011)) color_data = 12'b001100000111;
		if(({row_reg, col_reg}==14'b01011010101100)) color_data = 12'b010000000100;
		if(({row_reg, col_reg}==14'b01011010101101)) color_data = 12'b011000100100;
		if(({row_reg, col_reg}==14'b01011010101110)) color_data = 12'b011100100101;
		if(({row_reg, col_reg}==14'b01011010101111)) color_data = 12'b011000100101;
		if(({row_reg, col_reg}>=14'b01011010110000) && ({row_reg, col_reg}<14'b01011010110010)) color_data = 12'b010100110100;
		if(({row_reg, col_reg}>=14'b01011010110010) && ({row_reg, col_reg}<14'b01011010110100)) color_data = 12'b011000110100;
		if(({row_reg, col_reg}==14'b01011010110100)) color_data = 12'b010100100011;
		if(({row_reg, col_reg}==14'b01011010110101)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}==14'b01011010110110)) color_data = 12'b001100010001;
		if(({row_reg, col_reg}>=14'b01011010110111) && ({row_reg, col_reg}<14'b01011010111001)) color_data = 12'b001100010010;
		if(({row_reg, col_reg}==14'b01011010111001)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==14'b01011010111010)) color_data = 12'b101010001001;
		if(({row_reg, col_reg}==14'b01011010111011)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}>=14'b01011010111100) && ({row_reg, col_reg}<14'b01011010111110)) color_data = 12'b100101110111;
		if(({row_reg, col_reg}>=14'b01011010111110) && ({row_reg, col_reg}<14'b01011011000000)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==14'b01011011000000)) color_data = 12'b100101111000;
		if(({row_reg, col_reg}==14'b01011011000001)) color_data = 12'b101010001000;
		if(({row_reg, col_reg}==14'b01011011000010)) color_data = 12'b011001000100;
		if(({row_reg, col_reg}==14'b01011011000011)) color_data = 12'b001000000000;
		if(({row_reg, col_reg}==14'b01011011000100)) color_data = 12'b010100100011;
		if(({row_reg, col_reg}==14'b01011011000101)) color_data = 12'b101110001001;
		if(({row_reg, col_reg}>=14'b01011011000110) && ({row_reg, col_reg}<14'b01011011001010)) color_data = 12'b101001111001;
		if(({row_reg, col_reg}==14'b01011011001010)) color_data = 12'b101110001001;
		if(({row_reg, col_reg}==14'b01011011001011)) color_data = 12'b101001111000;
		if(({row_reg, col_reg}==14'b01011011001100)) color_data = 12'b101001111001;
		if(({row_reg, col_reg}==14'b01011011001101)) color_data = 12'b101110001001;
		if(({row_reg, col_reg}==14'b01011011001110)) color_data = 12'b101101111000;
		if(({row_reg, col_reg}==14'b01011011001111)) color_data = 12'b101110001001;
		if(({row_reg, col_reg}==14'b01011011010000)) color_data = 12'b100100100100;
		if(({row_reg, col_reg}==14'b01011011010001)) color_data = 12'b011100000010;
		if(({row_reg, col_reg}==14'b01011011010010)) color_data = 12'b100000010011;
		if(({row_reg, col_reg}==14'b01011011010011)) color_data = 12'b101000110101;
		if(({row_reg, col_reg}==14'b01011011010100)) color_data = 12'b101000110110;
		if(({row_reg, col_reg}==14'b01011011010101)) color_data = 12'b011100100111;
		if(({row_reg, col_reg}==14'b01011011010110)) color_data = 12'b010000001000;
		if(({row_reg, col_reg}==14'b01011011010111)) color_data = 12'b000100001011;
		if(({row_reg, col_reg}==14'b01011011011000)) color_data = 12'b000000001110;

		if(({row_reg, col_reg}>=14'b01011011011001) && ({row_reg, col_reg}<14'b01011100100111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==14'b01011100100111)) color_data = 12'b000000001110;
		if(({row_reg, col_reg}==14'b01011100101000)) color_data = 12'b000000001101;
		if(({row_reg, col_reg}==14'b01011100101001)) color_data = 12'b000100001011;
		if(({row_reg, col_reg}==14'b01011100101010)) color_data = 12'b001000001000;
		if(({row_reg, col_reg}==14'b01011100101011)) color_data = 12'b010000100110;
		if(({row_reg, col_reg}==14'b01011100101100)) color_data = 12'b010100010011;
		if(({row_reg, col_reg}==14'b01011100101101)) color_data = 12'b011000100100;
		if(({row_reg, col_reg}==14'b01011100101110)) color_data = 12'b011000110100;
		if(({row_reg, col_reg}==14'b01011100101111)) color_data = 12'b010100110100;
		if(({row_reg, col_reg}==14'b01011100110000)) color_data = 12'b010100110101;
		if(({row_reg, col_reg}==14'b01011100110001)) color_data = 12'b010100110100;
		if(({row_reg, col_reg}==14'b01011100110010)) color_data = 12'b010100100100;
		if(({row_reg, col_reg}>=14'b01011100110011) && ({row_reg, col_reg}<14'b01011100110101)) color_data = 12'b010000100011;
		if(({row_reg, col_reg}==14'b01011100110101)) color_data = 12'b001100010010;
		if(({row_reg, col_reg}==14'b01011100110110)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}>=14'b01011100110111) && ({row_reg, col_reg}<14'b01011100111001)) color_data = 12'b011001010101;
		if(({row_reg, col_reg}==14'b01011100111001)) color_data = 12'b100101111000;
		if(({row_reg, col_reg}==14'b01011100111010)) color_data = 12'b101010001001;
		if(({row_reg, col_reg}>=14'b01011100111011) && ({row_reg, col_reg}<14'b01011101000001)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==14'b01011101000001)) color_data = 12'b101010001000;
		if(({row_reg, col_reg}==14'b01011101000010)) color_data = 12'b011001000100;
		if(({row_reg, col_reg}==14'b01011101000011)) color_data = 12'b001000000000;
		if(({row_reg, col_reg}==14'b01011101000100)) color_data = 12'b010100110011;
		if(({row_reg, col_reg}==14'b01011101000101)) color_data = 12'b101010001001;
		if(({row_reg, col_reg}>=14'b01011101000110) && ({row_reg, col_reg}<14'b01011101001000)) color_data = 12'b100101111000;
		if(({row_reg, col_reg}>=14'b01011101001000) && ({row_reg, col_reg}<14'b01011101001011)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}>=14'b01011101001011) && ({row_reg, col_reg}<14'b01011101001101)) color_data = 12'b100101111000;
		if(({row_reg, col_reg}==14'b01011101001101)) color_data = 12'b100101110111;
		if(({row_reg, col_reg}>=14'b01011101001110) && ({row_reg, col_reg}<14'b01011101010000)) color_data = 12'b011101010101;
		if(({row_reg, col_reg}==14'b01011101010000)) color_data = 12'b011100110101;
		if(({row_reg, col_reg}==14'b01011101010001)) color_data = 12'b011000100011;
		if(({row_reg, col_reg}==14'b01011101010010)) color_data = 12'b011100100011;
		if(({row_reg, col_reg}==14'b01011101010011)) color_data = 12'b100000110100;
		if(({row_reg, col_reg}==14'b01011101010100)) color_data = 12'b100000100100;
		if(({row_reg, col_reg}==14'b01011101010101)) color_data = 12'b010100010101;
		if(({row_reg, col_reg}==14'b01011101010110)) color_data = 12'b001000000111;
		if(({row_reg, col_reg}==14'b01011101010111)) color_data = 12'b000100001011;
		if(({row_reg, col_reg}==14'b01011101011000)) color_data = 12'b000000001110;

		if(({row_reg, col_reg}>=14'b01011101011001) && ({row_reg, col_reg}<14'b01011110100110)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=14'b01011110100110) && ({row_reg, col_reg}<14'b01011110101000)) color_data = 12'b000000001110;
		if(({row_reg, col_reg}==14'b01011110101000)) color_data = 12'b000100001101;
		if(({row_reg, col_reg}==14'b01011110101001)) color_data = 12'b000000001010;
		if(({row_reg, col_reg}==14'b01011110101010)) color_data = 12'b001000000111;
		if(({row_reg, col_reg}==14'b01011110101011)) color_data = 12'b010100110110;
		if(({row_reg, col_reg}==14'b01011110101100)) color_data = 12'b011000110100;
		if(({row_reg, col_reg}==14'b01011110101101)) color_data = 12'b011000110011;
		if(({row_reg, col_reg}==14'b01011110101110)) color_data = 12'b011000110100;
		if(({row_reg, col_reg}>=14'b01011110101111) && ({row_reg, col_reg}<14'b01011110110010)) color_data = 12'b010100110101;
		if(({row_reg, col_reg}==14'b01011110110010)) color_data = 12'b010000100011;
		if(({row_reg, col_reg}>=14'b01011110110011) && ({row_reg, col_reg}<14'b01011110110101)) color_data = 12'b010000010011;
		if(({row_reg, col_reg}==14'b01011110110101)) color_data = 12'b001100010010;
		if(({row_reg, col_reg}==14'b01011110110110)) color_data = 12'b010000110011;
		if(({row_reg, col_reg}==14'b01011110110111)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==14'b01011110111000)) color_data = 12'b100110001001;
		if(({row_reg, col_reg}==14'b01011110111001)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==14'b01011110111010)) color_data = 12'b100001111000;
		if(({row_reg, col_reg}>=14'b01011110111011) && ({row_reg, col_reg}<14'b01011110111101)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==14'b01011110111101)) color_data = 12'b100001111000;
		if(({row_reg, col_reg}==14'b01011110111110)) color_data = 12'b100101111000;
		if(({row_reg, col_reg}>=14'b01011110111111) && ({row_reg, col_reg}<14'b01011111000010)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==14'b01011111000010)) color_data = 12'b011001000101;
		if(({row_reg, col_reg}==14'b01011111000011)) color_data = 12'b001000000000;
		if(({row_reg, col_reg}==14'b01011111000100)) color_data = 12'b010100110011;
		if(({row_reg, col_reg}==14'b01011111000101)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==14'b01011111000110)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}>=14'b01011111000111) && ({row_reg, col_reg}<14'b01011111001010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=14'b01011111001010) && ({row_reg, col_reg}<14'b01011111001100)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==14'b01011111001100)) color_data = 12'b101010001001;
		if(({row_reg, col_reg}==14'b01011111001101)) color_data = 12'b100101110111;
		if(({row_reg, col_reg}==14'b01011111001110)) color_data = 12'b010100110100;
		if(({row_reg, col_reg}==14'b01011111001111)) color_data = 12'b010100110011;
		if(({row_reg, col_reg}==14'b01011111010000)) color_data = 12'b010100110101;
		if(({row_reg, col_reg}==14'b01011111010001)) color_data = 12'b011000110101;
		if(({row_reg, col_reg}==14'b01011111010010)) color_data = 12'b011100110100;
		if(({row_reg, col_reg}==14'b01011111010011)) color_data = 12'b011100100011;
		if(({row_reg, col_reg}==14'b01011111010100)) color_data = 12'b011000100010;
		if(({row_reg, col_reg}==14'b01011111010101)) color_data = 12'b010000000011;
		if(({row_reg, col_reg}==14'b01011111010110)) color_data = 12'b000100000110;
		if(({row_reg, col_reg}==14'b01011111010111)) color_data = 12'b000100001010;
		if(({row_reg, col_reg}==14'b01011111011000)) color_data = 12'b000000001101;

		if(({row_reg, col_reg}>=14'b01011111011001) && ({row_reg, col_reg}<14'b01100000100011)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==14'b01100000100011)) color_data = 12'b000000001110;
		if(({row_reg, col_reg}==14'b01100000100100)) color_data = 12'b000100001101;
		if(({row_reg, col_reg}==14'b01100000100101)) color_data = 12'b000100001100;
		if(({row_reg, col_reg}==14'b01100000100110)) color_data = 12'b001000001011;
		if(({row_reg, col_reg}==14'b01100000100111)) color_data = 12'b001000001001;
		if(({row_reg, col_reg}==14'b01100000101000)) color_data = 12'b001000000111;
		if(({row_reg, col_reg}==14'b01100000101001)) color_data = 12'b001100100110;
		if(({row_reg, col_reg}==14'b01100000101010)) color_data = 12'b010000100101;
		if(({row_reg, col_reg}>=14'b01100000101011) && ({row_reg, col_reg}<14'b01100000101101)) color_data = 12'b010100110101;
		if(({row_reg, col_reg}==14'b01100000101101)) color_data = 12'b010100110100;
		if(({row_reg, col_reg}==14'b01100000101110)) color_data = 12'b010100100100;
		if(({row_reg, col_reg}>=14'b01100000101111) && ({row_reg, col_reg}<14'b01100000110001)) color_data = 12'b010100110100;
		if(({row_reg, col_reg}>=14'b01100000110001) && ({row_reg, col_reg}<14'b01100000110011)) color_data = 12'b010000100011;
		if(({row_reg, col_reg}==14'b01100000110011)) color_data = 12'b001100010010;
		if(({row_reg, col_reg}==14'b01100000110100)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==14'b01100000110101)) color_data = 12'b001100010010;
		if(({row_reg, col_reg}==14'b01100000110110)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}>=14'b01100000110111) && ({row_reg, col_reg}<14'b01100000111001)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}>=14'b01100000111001) && ({row_reg, col_reg}<14'b01100000111011)) color_data = 12'b100110001001;
		if(({row_reg, col_reg}>=14'b01100000111011) && ({row_reg, col_reg}<14'b01100000111101)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==14'b01100000111101)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==14'b01100000111110)) color_data = 12'b100110001001;
		if(({row_reg, col_reg}==14'b01100000111111)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==14'b01100001000000)) color_data = 12'b100110001001;
		if(({row_reg, col_reg}==14'b01100001000001)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==14'b01100001000010)) color_data = 12'b011001010101;
		if(({row_reg, col_reg}==14'b01100001000011)) color_data = 12'b001000000001;
		if(({row_reg, col_reg}==14'b01100001000100)) color_data = 12'b010101000100;
		if(({row_reg, col_reg}==14'b01100001000101)) color_data = 12'b101010001001;
		if(({row_reg, col_reg}==14'b01100001000110)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==14'b01100001000111)) color_data = 12'b100101111000;
		if(({row_reg, col_reg}>=14'b01100001001000) && ({row_reg, col_reg}<14'b01100001001101)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==14'b01100001001101)) color_data = 12'b100101111000;
		if(({row_reg, col_reg}>=14'b01100001001110) && ({row_reg, col_reg}<14'b01100001010000)) color_data = 12'b010100110100;
		if(({row_reg, col_reg}==14'b01100001010000)) color_data = 12'b011000110100;
		if(({row_reg, col_reg}>=14'b01100001010001) && ({row_reg, col_reg}<14'b01100001010100)) color_data = 12'b010100110100;
		if(({row_reg, col_reg}==14'b01100001010100)) color_data = 12'b010100110011;
		if(({row_reg, col_reg}==14'b01100001010101)) color_data = 12'b001100010100;
		if(({row_reg, col_reg}==14'b01100001010110)) color_data = 12'b000000000110;
		if(({row_reg, col_reg}==14'b01100001010111)) color_data = 12'b000000001011;
		if(({row_reg, col_reg}==14'b01100001011000)) color_data = 12'b000000001110;

		if(({row_reg, col_reg}>=14'b01100001011001) && ({row_reg, col_reg}<14'b01100010100010)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==14'b01100010100010)) color_data = 12'b000000001110;
		if(({row_reg, col_reg}==14'b01100010100011)) color_data = 12'b000100001100;
		if(({row_reg, col_reg}==14'b01100010100100)) color_data = 12'b000100001010;
		if(({row_reg, col_reg}==14'b01100010100101)) color_data = 12'b001000001001;
		if(({row_reg, col_reg}==14'b01100010100110)) color_data = 12'b001100011001;
		if(({row_reg, col_reg}==14'b01100010100111)) color_data = 12'b001100000111;
		if(({row_reg, col_reg}==14'b01100010101000)) color_data = 12'b001100010110;
		if(({row_reg, col_reg}==14'b01100010101001)) color_data = 12'b010000100110;
		if(({row_reg, col_reg}>=14'b01100010101010) && ({row_reg, col_reg}<14'b01100010101100)) color_data = 12'b010100110101;
		if(({row_reg, col_reg}==14'b01100010101100)) color_data = 12'b011000110100;
		if(({row_reg, col_reg}==14'b01100010101101)) color_data = 12'b010100100011;
		if(({row_reg, col_reg}>=14'b01100010101110) && ({row_reg, col_reg}<14'b01100010110100)) color_data = 12'b001100010010;
		if(({row_reg, col_reg}>=14'b01100010110100) && ({row_reg, col_reg}<14'b01100010110110)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==14'b01100010110110)) color_data = 12'b010000100011;
		if(({row_reg, col_reg}==14'b01100010110111)) color_data = 12'b100101111000;
		if(({row_reg, col_reg}==14'b01100010111000)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==14'b01100010111001)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}>=14'b01100010111010) && ({row_reg, col_reg}<14'b01100010111100)) color_data = 12'b110010111011;
		if(({row_reg, col_reg}>=14'b01100010111100) && ({row_reg, col_reg}<14'b01100010111111)) color_data = 12'b110010101011;
		if(({row_reg, col_reg}==14'b01100010111111)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}>=14'b01100011000000) && ({row_reg, col_reg}<14'b01100011000010)) color_data = 12'b110010111011;
		if(({row_reg, col_reg}==14'b01100011000010)) color_data = 12'b011001010101;
		if(({row_reg, col_reg}==14'b01100011000011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==14'b01100011000100)) color_data = 12'b010101000100;
		if(({row_reg, col_reg}>=14'b01100011000101) && ({row_reg, col_reg}<14'b01100011000111)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==14'b01100011000111)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}>=14'b01100011001000) && ({row_reg, col_reg}<14'b01100011001101)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==14'b01100011001101)) color_data = 12'b100101111000;
		if(({row_reg, col_reg}>=14'b01100011001110) && ({row_reg, col_reg}<14'b01100011010101)) color_data = 12'b010100110100;
		if(({row_reg, col_reg}==14'b01100011010101)) color_data = 12'b001100010100;
		if(({row_reg, col_reg}==14'b01100011010110)) color_data = 12'b000000000110;
		if(({row_reg, col_reg}==14'b01100011010111)) color_data = 12'b000000001010;
		if(({row_reg, col_reg}==14'b01100011011000)) color_data = 12'b000000001110;

		if(({row_reg, col_reg}>=14'b01100011011001) && ({row_reg, col_reg}<14'b01100100100001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==14'b01100100100001)) color_data = 12'b000000001110;
		if(({row_reg, col_reg}==14'b01100100100010)) color_data = 12'b000100001100;
		if(({row_reg, col_reg}==14'b01100100100011)) color_data = 12'b001000001010;
		if(({row_reg, col_reg}==14'b01100100100100)) color_data = 12'b001100011000;
		if(({row_reg, col_reg}==14'b01100100100101)) color_data = 12'b010100101000;
		if(({row_reg, col_reg}==14'b01100100100110)) color_data = 12'b011000110111;
		if(({row_reg, col_reg}==14'b01100100100111)) color_data = 12'b010100110110;
		if(({row_reg, col_reg}>=14'b01100100101000) && ({row_reg, col_reg}<14'b01100100101010)) color_data = 12'b010100110101;
		if(({row_reg, col_reg}>=14'b01100100101010) && ({row_reg, col_reg}<14'b01100100101100)) color_data = 12'b010100110100;
		if(({row_reg, col_reg}==14'b01100100101100)) color_data = 12'b011000110100;
		if(({row_reg, col_reg}==14'b01100100101101)) color_data = 12'b010100100011;
		if(({row_reg, col_reg}==14'b01100100101110)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}>=14'b01100100101111) && ({row_reg, col_reg}<14'b01100100110010)) color_data = 12'b001100010010;
		if(({row_reg, col_reg}>=14'b01100100110010) && ({row_reg, col_reg}<14'b01100100110100)) color_data = 12'b010000100011;
		if(({row_reg, col_reg}==14'b01100100110100)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==14'b01100100110101)) color_data = 12'b001100010010;
		if(({row_reg, col_reg}==14'b01100100110110)) color_data = 12'b010000100011;
		if(({row_reg, col_reg}>=14'b01100100110111) && ({row_reg, col_reg}<14'b01100100111001)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==14'b01100100111001)) color_data = 12'b101110011010;
		if(({row_reg, col_reg}>=14'b01100100111010) && ({row_reg, col_reg}<14'b01100100111100)) color_data = 12'b101110101011;
		if(({row_reg, col_reg}>=14'b01100100111100) && ({row_reg, col_reg}<14'b01100100111110)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==14'b01100100111110)) color_data = 12'b110010111011;
		if(({row_reg, col_reg}>=14'b01100100111111) && ({row_reg, col_reg}<14'b01100101000001)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==14'b01100101000001)) color_data = 12'b110010111011;
		if(({row_reg, col_reg}==14'b01100101000010)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==14'b01100101000011)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==14'b01100101000100)) color_data = 12'b011001000101;
		if(({row_reg, col_reg}==14'b01100101000101)) color_data = 12'b110010111011;
		if(({row_reg, col_reg}==14'b01100101000110)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==14'b01100101000111)) color_data = 12'b100101111000;
		if(({row_reg, col_reg}>=14'b01100101001000) && ({row_reg, col_reg}<14'b01100101001101)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==14'b01100101001101)) color_data = 12'b100101111000;
		if(({row_reg, col_reg}>=14'b01100101001110) && ({row_reg, col_reg}<14'b01100101010001)) color_data = 12'b010100110100;
		if(({row_reg, col_reg}==14'b01100101010001)) color_data = 12'b011000110100;
		if(({row_reg, col_reg}==14'b01100101010010)) color_data = 12'b010100110100;
		if(({row_reg, col_reg}==14'b01100101010011)) color_data = 12'b010100100011;
		if(({row_reg, col_reg}==14'b01100101010100)) color_data = 12'b010100110100;
		if(({row_reg, col_reg}==14'b01100101010101)) color_data = 12'b001100010100;
		if(({row_reg, col_reg}==14'b01100101010110)) color_data = 12'b000100000110;
		if(({row_reg, col_reg}==14'b01100101010111)) color_data = 12'b000000001010;
		if(({row_reg, col_reg}==14'b01100101011000)) color_data = 12'b000000001101;

		if(({row_reg, col_reg}>=14'b01100101011001) && ({row_reg, col_reg}<14'b01100110100000)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==14'b01100110100000)) color_data = 12'b000000001110;
		if(({row_reg, col_reg}==14'b01100110100001)) color_data = 12'b001000001101;
		if(({row_reg, col_reg}==14'b01100110100010)) color_data = 12'b001100001010;
		if(({row_reg, col_reg}==14'b01100110100011)) color_data = 12'b010100011000;
		if(({row_reg, col_reg}==14'b01100110100100)) color_data = 12'b011000100110;
		if(({row_reg, col_reg}==14'b01100110100101)) color_data = 12'b011000110101;
		if(({row_reg, col_reg}==14'b01100110100110)) color_data = 12'b011000110100;
		if(({row_reg, col_reg}==14'b01100110100111)) color_data = 12'b010100110011;
		if(({row_reg, col_reg}==14'b01100110101000)) color_data = 12'b011000110100;
		if(({row_reg, col_reg}>=14'b01100110101001) && ({row_reg, col_reg}<14'b01100110101100)) color_data = 12'b010100110100;
		if(({row_reg, col_reg}==14'b01100110101100)) color_data = 12'b011000110100;
		if(({row_reg, col_reg}>=14'b01100110101101) && ({row_reg, col_reg}<14'b01100110110000)) color_data = 12'b010100110100;
		if(({row_reg, col_reg}==14'b01100110110000)) color_data = 12'b010000010010;
		if(({row_reg, col_reg}==14'b01100110110001)) color_data = 12'b001100010010;
		if(({row_reg, col_reg}==14'b01100110110010)) color_data = 12'b010000100011;
		if(({row_reg, col_reg}==14'b01100110110011)) color_data = 12'b010100110100;
		if(({row_reg, col_reg}==14'b01100110110100)) color_data = 12'b010000110011;
		if(({row_reg, col_reg}==14'b01100110110101)) color_data = 12'b001100010010;
		if(({row_reg, col_reg}==14'b01100110110110)) color_data = 12'b010000110011;
		if(({row_reg, col_reg}>=14'b01100110110111) && ({row_reg, col_reg}<14'b01100110111011)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==14'b01100110111011)) color_data = 12'b110010101011;
		if(({row_reg, col_reg}>=14'b01100110111100) && ({row_reg, col_reg}<14'b01100110111110)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==14'b01100110111110)) color_data = 12'b110010111011;
		if(({row_reg, col_reg}>=14'b01100110111111) && ({row_reg, col_reg}<14'b01100111000001)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==14'b01100111000001)) color_data = 12'b110010111011;
		if(({row_reg, col_reg}==14'b01100111000010)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==14'b01100111000011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}==14'b01100111000100)) color_data = 12'b010100110100;
		if(({row_reg, col_reg}>=14'b01100111000101) && ({row_reg, col_reg}<14'b01100111000111)) color_data = 12'b110010111011;
		if(({row_reg, col_reg}>=14'b01100111000111) && ({row_reg, col_reg}<14'b01100111001011)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==14'b01100111001011)) color_data = 12'b100101111000;
		if(({row_reg, col_reg}==14'b01100111001100)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==14'b01100111001101)) color_data = 12'b100101111000;
		if(({row_reg, col_reg}>=14'b01100111001110) && ({row_reg, col_reg}<14'b01100111010001)) color_data = 12'b010100110100;
		if(({row_reg, col_reg}==14'b01100111010001)) color_data = 12'b011000110100;
		if(({row_reg, col_reg}==14'b01100111010010)) color_data = 12'b010000100011;
		if(({row_reg, col_reg}==14'b01100111010011)) color_data = 12'b001100010010;
		if(({row_reg, col_reg}==14'b01100111010100)) color_data = 12'b010000010011;
		if(({row_reg, col_reg}==14'b01100111010101)) color_data = 12'b001000010011;
		if(({row_reg, col_reg}==14'b01100111010110)) color_data = 12'b000100000101;
		if(({row_reg, col_reg}==14'b01100111010111)) color_data = 12'b000000001001;
		if(({row_reg, col_reg}==14'b01100111011000)) color_data = 12'b000000001100;
		if(({row_reg, col_reg}==14'b01100111011001)) color_data = 12'b000000001110;

		if(({row_reg, col_reg}>=14'b01100111011010) && ({row_reg, col_reg}<14'b01101000100000)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==14'b01101000100000)) color_data = 12'b000100001100;
		if(({row_reg, col_reg}==14'b01101000100001)) color_data = 12'b001100001011;
		if(({row_reg, col_reg}==14'b01101000100010)) color_data = 12'b010100011001;
		if(({row_reg, col_reg}==14'b01101000100011)) color_data = 12'b100000100111;
		if(({row_reg, col_reg}==14'b01101000100100)) color_data = 12'b100000110101;
		if(({row_reg, col_reg}==14'b01101000100101)) color_data = 12'b011100100011;
		if(({row_reg, col_reg}>=14'b01101000100110) && ({row_reg, col_reg}<14'b01101000101000)) color_data = 12'b011000110011;
		if(({row_reg, col_reg}==14'b01101000101000)) color_data = 12'b010100110011;
		if(({row_reg, col_reg}>=14'b01101000101001) && ({row_reg, col_reg}<14'b01101000101100)) color_data = 12'b010100110100;
		if(({row_reg, col_reg}==14'b01101000101100)) color_data = 12'b011000110100;
		if(({row_reg, col_reg}>=14'b01101000101101) && ({row_reg, col_reg}<14'b01101000110000)) color_data = 12'b010100110100;
		if(({row_reg, col_reg}>=14'b01101000110000) && ({row_reg, col_reg}<14'b01101000110010)) color_data = 12'b010000010010;
		if(({row_reg, col_reg}==14'b01101000110010)) color_data = 12'b010100100011;
		if(({row_reg, col_reg}>=14'b01101000110011) && ({row_reg, col_reg}<14'b01101000110101)) color_data = 12'b010100110100;
		if(({row_reg, col_reg}==14'b01101000110101)) color_data = 12'b001100010010;
		if(({row_reg, col_reg}==14'b01101000110110)) color_data = 12'b010000100011;
		if(({row_reg, col_reg}>=14'b01101000110111) && ({row_reg, col_reg}<14'b01101000111010)) color_data = 12'b110010101011;
		if(({row_reg, col_reg}==14'b01101000111010)) color_data = 12'b101110101011;
		if(({row_reg, col_reg}>=14'b01101000111011) && ({row_reg, col_reg}<14'b01101000111101)) color_data = 12'b110010111011;
		if(({row_reg, col_reg}==14'b01101000111101)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}>=14'b01101000111110) && ({row_reg, col_reg}<14'b01101001000000)) color_data = 12'b101110101011;
		if(({row_reg, col_reg}==14'b01101001000000)) color_data = 12'b110010111011;
		if(({row_reg, col_reg}==14'b01101001000001)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==14'b01101001000010)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==14'b01101001000011)) color_data = 12'b001000000001;
		if(({row_reg, col_reg}==14'b01101001000100)) color_data = 12'b010101000100;
		if(({row_reg, col_reg}>=14'b01101001000101) && ({row_reg, col_reg}<14'b01101001000111)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}>=14'b01101001000111) && ({row_reg, col_reg}<14'b01101001001011)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==14'b01101001001011)) color_data = 12'b100101111000;
		if(({row_reg, col_reg}==14'b01101001001100)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==14'b01101001001101)) color_data = 12'b100101111000;
		if(({row_reg, col_reg}>=14'b01101001001110) && ({row_reg, col_reg}<14'b01101001010010)) color_data = 12'b010100110100;
		if(({row_reg, col_reg}==14'b01101001010010)) color_data = 12'b010000100011;
		if(({row_reg, col_reg}>=14'b01101001010011) && ({row_reg, col_reg}<14'b01101001010101)) color_data = 12'b001100010010;
		if(({row_reg, col_reg}==14'b01101001010101)) color_data = 12'b001000000011;
		if(({row_reg, col_reg}==14'b01101001010110)) color_data = 12'b000100000100;
		if(({row_reg, col_reg}==14'b01101001010111)) color_data = 12'b000100001000;
		if(({row_reg, col_reg}==14'b01101001011000)) color_data = 12'b000000001011;
		if(({row_reg, col_reg}==14'b01101001011001)) color_data = 12'b000000001101;

		if(({row_reg, col_reg}>=14'b01101001011010) && ({row_reg, col_reg}<14'b01101010011110)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=14'b01101010011110) && ({row_reg, col_reg}<14'b01101010100000)) color_data = 12'b000000001110;
		if(({row_reg, col_reg}==14'b01101010100000)) color_data = 12'b010000001001;
		if(({row_reg, col_reg}==14'b01101010100001)) color_data = 12'b011000011001;
		if(({row_reg, col_reg}==14'b01101010100010)) color_data = 12'b100000101000;
		if(({row_reg, col_reg}==14'b01101010100011)) color_data = 12'b101000110110;
		if(({row_reg, col_reg}==14'b01101010100100)) color_data = 12'b100000100011;
		if(({row_reg, col_reg}==14'b01101010100101)) color_data = 12'b011000010001;
		if(({row_reg, col_reg}==14'b01101010100110)) color_data = 12'b010100100001;
		if(({row_reg, col_reg}==14'b01101010100111)) color_data = 12'b011000110011;
		if(({row_reg, col_reg}>=14'b01101010101000) && ({row_reg, col_reg}<14'b01101010101010)) color_data = 12'b010100110100;
		if(({row_reg, col_reg}==14'b01101010101010)) color_data = 12'b010100110101;
		if(({row_reg, col_reg}>=14'b01101010101011) && ({row_reg, col_reg}<14'b01101010110000)) color_data = 12'b010100110100;
		if(({row_reg, col_reg}>=14'b01101010110000) && ({row_reg, col_reg}<14'b01101010110010)) color_data = 12'b010100100011;
		if(({row_reg, col_reg}>=14'b01101010110010) && ({row_reg, col_reg}<14'b01101010110101)) color_data = 12'b010000100011;
		if(({row_reg, col_reg}==14'b01101010110101)) color_data = 12'b001100010010;
		if(({row_reg, col_reg}==14'b01101010110110)) color_data = 12'b010000100011;
		if(({row_reg, col_reg}>=14'b01101010110111) && ({row_reg, col_reg}<14'b01101010111001)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}>=14'b01101010111001) && ({row_reg, col_reg}<14'b01101010111011)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==14'b01101010111011)) color_data = 12'b101110101011;
		if(({row_reg, col_reg}>=14'b01101010111100) && ({row_reg, col_reg}<14'b01101010111110)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==14'b01101010111110)) color_data = 12'b101110101011;
		if(({row_reg, col_reg}==14'b01101010111111)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==14'b01101011000000)) color_data = 12'b011001010101;
		if(({row_reg, col_reg}==14'b01101011000001)) color_data = 12'b010101000100;
		if(({row_reg, col_reg}==14'b01101011000010)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==14'b01101011000011)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==14'b01101011000100)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==14'b01101011000101)) color_data = 12'b110010111011;
		if(({row_reg, col_reg}==14'b01101011000110)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}>=14'b01101011000111) && ({row_reg, col_reg}<14'b01101011001011)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==14'b01101011001011)) color_data = 12'b100101111000;
		if(({row_reg, col_reg}==14'b01101011001100)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==14'b01101011001101)) color_data = 12'b100101111000;
		if(({row_reg, col_reg}>=14'b01101011001110) && ({row_reg, col_reg}<14'b01101011010011)) color_data = 12'b010100110100;
		if(({row_reg, col_reg}==14'b01101011010011)) color_data = 12'b010100100011;
		if(({row_reg, col_reg}==14'b01101011010100)) color_data = 12'b010000100011;
		if(({row_reg, col_reg}==14'b01101011010101)) color_data = 12'b001100010011;
		if(({row_reg, col_reg}==14'b01101011010110)) color_data = 12'b001000000011;
		if(({row_reg, col_reg}==14'b01101011010111)) color_data = 12'b000100000110;
		if(({row_reg, col_reg}==14'b01101011011000)) color_data = 12'b000000001001;
		if(({row_reg, col_reg}==14'b01101011011001)) color_data = 12'b000000001100;
		if(({row_reg, col_reg}==14'b01101011011010)) color_data = 12'b000000001110;

		if(({row_reg, col_reg}>=14'b01101011011011) && ({row_reg, col_reg}<14'b01101100011101)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==14'b01101100011101)) color_data = 12'b000000001110;
		if(({row_reg, col_reg}==14'b01101100011110)) color_data = 12'b000100001100;
		if(({row_reg, col_reg}==14'b01101100011111)) color_data = 12'b001000001100;
		if(({row_reg, col_reg}==14'b01101100100000)) color_data = 12'b011000000110;
		if(({row_reg, col_reg}==14'b01101100100001)) color_data = 12'b100000010110;
		if(({row_reg, col_reg}==14'b01101100100010)) color_data = 12'b101000100110;
		if(({row_reg, col_reg}==14'b01101100100011)) color_data = 12'b101100100101;
		if(({row_reg, col_reg}==14'b01101100100100)) color_data = 12'b100000010010;
		if(({row_reg, col_reg}==14'b01101100100101)) color_data = 12'b010100000001;
		if(({row_reg, col_reg}==14'b01101100100110)) color_data = 12'b010100010010;
		if(({row_reg, col_reg}==14'b01101100100111)) color_data = 12'b011000110100;
		if(({row_reg, col_reg}>=14'b01101100101000) && ({row_reg, col_reg}<14'b01101100110010)) color_data = 12'b010100110100;
		if(({row_reg, col_reg}==14'b01101100110010)) color_data = 12'b010000100011;
		if(({row_reg, col_reg}>=14'b01101100110011) && ({row_reg, col_reg}<14'b01101100110110)) color_data = 12'b001100010010;
		if(({row_reg, col_reg}==14'b01101100110110)) color_data = 12'b010000100011;
		if(({row_reg, col_reg}==14'b01101100110111)) color_data = 12'b100101111000;
		if(({row_reg, col_reg}==14'b01101100111000)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==14'b01101100111001)) color_data = 12'b110010101011;
		if(({row_reg, col_reg}==14'b01101100111010)) color_data = 12'b110010111011;
		if(({row_reg, col_reg}==14'b01101100111011)) color_data = 12'b101110101011;
		if(({row_reg, col_reg}==14'b01101100111100)) color_data = 12'b110010101011;
		if(({row_reg, col_reg}==14'b01101100111101)) color_data = 12'b101110101011;
		if(({row_reg, col_reg}>=14'b01101100111110) && ({row_reg, col_reg}<14'b01101101000000)) color_data = 12'b110010111011;
		if(({row_reg, col_reg}==14'b01101101000000)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==14'b01101101000001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==14'b01101101000010)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==14'b01101101000011)) color_data = 12'b110110111100;
		if(({row_reg, col_reg}==14'b01101101000100)) color_data = 12'b110010111011;
		if(({row_reg, col_reg}==14'b01101101000101)) color_data = 12'b110010101011;
		if(({row_reg, col_reg}==14'b01101101000110)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==14'b01101101000111)) color_data = 12'b100110001001;
		if(({row_reg, col_reg}>=14'b01101101001000) && ({row_reg, col_reg}<14'b01101101001011)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==14'b01101101001011)) color_data = 12'b100101111000;
		if(({row_reg, col_reg}==14'b01101101001100)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==14'b01101101001101)) color_data = 12'b100101111000;
		if(({row_reg, col_reg}>=14'b01101101001110) && ({row_reg, col_reg}<14'b01101101010100)) color_data = 12'b010100110100;
		if(({row_reg, col_reg}==14'b01101101010100)) color_data = 12'b010100100011;
		if(({row_reg, col_reg}==14'b01101101010101)) color_data = 12'b001100010010;
		if(({row_reg, col_reg}==14'b01101101010110)) color_data = 12'b001000010011;
		if(({row_reg, col_reg}==14'b01101101010111)) color_data = 12'b000100000101;
		if(({row_reg, col_reg}==14'b01101101011000)) color_data = 12'b000000000111;
		if(({row_reg, col_reg}==14'b01101101011001)) color_data = 12'b000000001011;
		if(({row_reg, col_reg}==14'b01101101011010)) color_data = 12'b000000001110;

		if(({row_reg, col_reg}>=14'b01101101011011) && ({row_reg, col_reg}<14'b01101110011100)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==14'b01101110011100)) color_data = 12'b000000001110;
		if(({row_reg, col_reg}==14'b01101110011101)) color_data = 12'b000100001100;
		if(({row_reg, col_reg}==14'b01101110011110)) color_data = 12'b001100001010;
		if(({row_reg, col_reg}==14'b01101110011111)) color_data = 12'b010000001001;
		if(({row_reg, col_reg}==14'b01101110100000)) color_data = 12'b100100010100;
		if(({row_reg, col_reg}==14'b01101110100001)) color_data = 12'b101000100101;
		if(({row_reg, col_reg}==14'b01101110100010)) color_data = 12'b101100100101;
		if(({row_reg, col_reg}==14'b01101110100011)) color_data = 12'b101100100100;
		if(({row_reg, col_reg}==14'b01101110100100)) color_data = 12'b100000010011;
		if(({row_reg, col_reg}==14'b01101110100101)) color_data = 12'b010100000001;
		if(({row_reg, col_reg}==14'b01101110100110)) color_data = 12'b010000010010;
		if(({row_reg, col_reg}>=14'b01101110100111) && ({row_reg, col_reg}<14'b01101110101101)) color_data = 12'b010100110100;
		if(({row_reg, col_reg}==14'b01101110101101)) color_data = 12'b011000110100;
		if(({row_reg, col_reg}==14'b01101110101110)) color_data = 12'b010100110100;
		if(({row_reg, col_reg}==14'b01101110101111)) color_data = 12'b010100110011;
		if(({row_reg, col_reg}==14'b01101110110000)) color_data = 12'b011000110100;
		if(({row_reg, col_reg}>=14'b01101110110001) && ({row_reg, col_reg}<14'b01101110110011)) color_data = 12'b010100110100;
		if(({row_reg, col_reg}>=14'b01101110110011) && ({row_reg, col_reg}<14'b01101110110111)) color_data = 12'b010000100011;
		if(({row_reg, col_reg}==14'b01101110110111)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==14'b01101110111000)) color_data = 12'b011101010110;
		if(({row_reg, col_reg}==14'b01101110111001)) color_data = 12'b101010001001;
		if(({row_reg, col_reg}==14'b01101110111010)) color_data = 12'b101110011010;
		if(({row_reg, col_reg}==14'b01101110111011)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==14'b01101110111100)) color_data = 12'b101110101011;
		if(({row_reg, col_reg}>=14'b01101110111101) && ({row_reg, col_reg}<14'b01101110111111)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==14'b01101110111111)) color_data = 12'b101110101011;
		if(({row_reg, col_reg}==14'b01101111000000)) color_data = 12'b010100110011;
		if(({row_reg, col_reg}==14'b01101111000001)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==14'b01101111000010)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==14'b01101111000011)) color_data = 12'b110010111011;
		if(({row_reg, col_reg}==14'b01101111000100)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}>=14'b01101111000101) && ({row_reg, col_reg}<14'b01101111000111)) color_data = 12'b101110011010;
		if(({row_reg, col_reg}>=14'b01101111000111) && ({row_reg, col_reg}<14'b01101111001011)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==14'b01101111001011)) color_data = 12'b100101111000;
		if(({row_reg, col_reg}==14'b01101111001100)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==14'b01101111001101)) color_data = 12'b100101111000;
		if(({row_reg, col_reg}>=14'b01101111001110) && ({row_reg, col_reg}<14'b01101111010100)) color_data = 12'b010100110100;
		if(({row_reg, col_reg}==14'b01101111010100)) color_data = 12'b010100110011;
		if(({row_reg, col_reg}==14'b01101111010101)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}==14'b01101111010110)) color_data = 12'b001100100011;
		if(({row_reg, col_reg}==14'b01101111010111)) color_data = 12'b001000010100;
		if(({row_reg, col_reg}==14'b01101111011000)) color_data = 12'b000000000110;
		if(({row_reg, col_reg}==14'b01101111011001)) color_data = 12'b000000001010;
		if(({row_reg, col_reg}==14'b01101111011010)) color_data = 12'b000000001101;

		if(({row_reg, col_reg}>=14'b01101111011011) && ({row_reg, col_reg}<14'b01110000011011)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==14'b01110000011011)) color_data = 12'b000000001110;
		if(({row_reg, col_reg}==14'b01110000011100)) color_data = 12'b000100001100;
		if(({row_reg, col_reg}==14'b01110000011101)) color_data = 12'b001100001001;
		if(({row_reg, col_reg}==14'b01110000011110)) color_data = 12'b011000001000;
		if(({row_reg, col_reg}==14'b01110000011111)) color_data = 12'b100000010111;
		if(({row_reg, col_reg}>=14'b01110000100000) && ({row_reg, col_reg}<14'b01110000100100)) color_data = 12'b101100100100;
		if(({row_reg, col_reg}==14'b01110000100100)) color_data = 12'b100000100011;
		if(({row_reg, col_reg}==14'b01110000100101)) color_data = 12'b010100000010;
		if(({row_reg, col_reg}>=14'b01110000100110) && ({row_reg, col_reg}<14'b01110000101001)) color_data = 12'b001100010010;
		if(({row_reg, col_reg}>=14'b01110000101001) && ({row_reg, col_reg}<14'b01110000101111)) color_data = 12'b010100110100;
		if(({row_reg, col_reg}==14'b01110000101111)) color_data = 12'b011000110100;
		if(({row_reg, col_reg}>=14'b01110000110000) && ({row_reg, col_reg}<14'b01110000110011)) color_data = 12'b010100110100;
		if(({row_reg, col_reg}==14'b01110000110011)) color_data = 12'b011000110100;
		if(({row_reg, col_reg}>=14'b01110000110100) && ({row_reg, col_reg}<14'b01110000110111)) color_data = 12'b010100110100;
		if(({row_reg, col_reg}==14'b01110000110111)) color_data = 12'b001100010010;
		if(({row_reg, col_reg}==14'b01110000111000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==14'b01110000111001)) color_data = 12'b100001100111;
		if(({row_reg, col_reg}==14'b01110000111010)) color_data = 12'b100101111000;
		if(({row_reg, col_reg}==14'b01110000111011)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==14'b01110000111100)) color_data = 12'b110010111011;
		if(({row_reg, col_reg}==14'b01110000111101)) color_data = 12'b110010101011;
		if(({row_reg, col_reg}==14'b01110000111110)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==14'b01110000111111)) color_data = 12'b101110101011;
		if(({row_reg, col_reg}==14'b01110001000000)) color_data = 12'b010000110011;
		if(({row_reg, col_reg}==14'b01110001000001)) color_data = 12'b001000000000;
		if(({row_reg, col_reg}==14'b01110001000010)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==14'b01110001000011)) color_data = 12'b110010111011;
		if(({row_reg, col_reg}==14'b01110001000100)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}>=14'b01110001000101) && ({row_reg, col_reg}<14'b01110001001001)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==14'b01110001001001)) color_data = 12'b100110001001;
		if(({row_reg, col_reg}==14'b01110001001010)) color_data = 12'b100101111000;
		if(({row_reg, col_reg}==14'b01110001001011)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==14'b01110001001100)) color_data = 12'b101010001001;
		if(({row_reg, col_reg}==14'b01110001001101)) color_data = 12'b101010001000;
		if(({row_reg, col_reg}>=14'b01110001001110) && ({row_reg, col_reg}<14'b01110001010001)) color_data = 12'b010100110100;
		if(({row_reg, col_reg}==14'b01110001010001)) color_data = 12'b010101000100;
		if(({row_reg, col_reg}>=14'b01110001010010) && ({row_reg, col_reg}<14'b01110001010101)) color_data = 12'b010100110100;
		if(({row_reg, col_reg}==14'b01110001010101)) color_data = 12'b010100110011;
		if(({row_reg, col_reg}==14'b01110001010110)) color_data = 12'b010100110100;
		if(({row_reg, col_reg}==14'b01110001010111)) color_data = 12'b001100100100;
		if(({row_reg, col_reg}==14'b01110001011000)) color_data = 12'b000000000101;
		if(({row_reg, col_reg}==14'b01110001011001)) color_data = 12'b000000001001;
		if(({row_reg, col_reg}==14'b01110001011010)) color_data = 12'b000000001101;

		if(({row_reg, col_reg}>=14'b01110001011011) && ({row_reg, col_reg}<14'b01110010011000)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==14'b01110010011000)) color_data = 12'b000000001110;
		if(({row_reg, col_reg}==14'b01110010011001)) color_data = 12'b000000001101;
		if(({row_reg, col_reg}==14'b01110010011010)) color_data = 12'b000100001100;
		if(({row_reg, col_reg}==14'b01110010011011)) color_data = 12'b001000001011;
		if(({row_reg, col_reg}==14'b01110010011100)) color_data = 12'b001100001001;
		if(({row_reg, col_reg}==14'b01110010011101)) color_data = 12'b011000001000;
		if(({row_reg, col_reg}==14'b01110010011110)) color_data = 12'b100000000110;
		if(({row_reg, col_reg}==14'b01110010011111)) color_data = 12'b101100010110;
		if(({row_reg, col_reg}>=14'b01110010100000) && ({row_reg, col_reg}<14'b01110010100011)) color_data = 12'b101100100100;
		if(({row_reg, col_reg}==14'b01110010100011)) color_data = 12'b101000100100;
		if(({row_reg, col_reg}==14'b01110010100100)) color_data = 12'b100000010011;
		if(({row_reg, col_reg}==14'b01110010100101)) color_data = 12'b010000010010;
		if(({row_reg, col_reg}==14'b01110010100110)) color_data = 12'b001100010011;
		if(({row_reg, col_reg}==14'b01110010100111)) color_data = 12'b001100010010;
		if(({row_reg, col_reg}==14'b01110010101000)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}>=14'b01110010101001) && ({row_reg, col_reg}<14'b01110010101011)) color_data = 12'b010100110011;
		if(({row_reg, col_reg}>=14'b01110010101011) && ({row_reg, col_reg}<14'b01110010110000)) color_data = 12'b010100110100;
		if(({row_reg, col_reg}==14'b01110010110000)) color_data = 12'b011000110101;
		if(({row_reg, col_reg}==14'b01110010110001)) color_data = 12'b011000110100;
		if(({row_reg, col_reg}>=14'b01110010110010) && ({row_reg, col_reg}<14'b01110010110111)) color_data = 12'b010100110100;
		if(({row_reg, col_reg}==14'b01110010110111)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}==14'b01110010111000)) color_data = 12'b001100010010;
		if(({row_reg, col_reg}==14'b01110010111001)) color_data = 12'b100001100111;
		if(({row_reg, col_reg}==14'b01110010111010)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==14'b01110010111011)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==14'b01110010111100)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==14'b01110010111101)) color_data = 12'b101110101011;
		if(({row_reg, col_reg}==14'b01110010111110)) color_data = 12'b110010111011;
		if(({row_reg, col_reg}==14'b01110010111111)) color_data = 12'b101110101011;
		if(({row_reg, col_reg}==14'b01110011000000)) color_data = 12'b010000110011;
		if(({row_reg, col_reg}==14'b01110011000001)) color_data = 12'b001000000000;
		if(({row_reg, col_reg}==14'b01110011000010)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==14'b01110011000011)) color_data = 12'b110010111011;
		if(({row_reg, col_reg}==14'b01110011000100)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}>=14'b01110011000101) && ({row_reg, col_reg}<14'b01110011001010)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}>=14'b01110011001010) && ({row_reg, col_reg}<14'b01110011001100)) color_data = 12'b100101111000;
		if(({row_reg, col_reg}>=14'b01110011001100) && ({row_reg, col_reg}<14'b01110011001110)) color_data = 12'b100001100111;
		if(({row_reg, col_reg}>=14'b01110011001110) && ({row_reg, col_reg}<14'b01110011010101)) color_data = 12'b010100110100;
		if(({row_reg, col_reg}==14'b01110011010101)) color_data = 12'b010100110011;
		if(({row_reg, col_reg}==14'b01110011010110)) color_data = 12'b010100110100;
		if(({row_reg, col_reg}==14'b01110011010111)) color_data = 12'b001100100011;
		if(({row_reg, col_reg}==14'b01110011011000)) color_data = 12'b000000000100;
		if(({row_reg, col_reg}==14'b01110011011001)) color_data = 12'b000000001001;
		if(({row_reg, col_reg}==14'b01110011011010)) color_data = 12'b000000001101;

		if(({row_reg, col_reg}>=14'b01110011011011) && ({row_reg, col_reg}<14'b01110100010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==14'b01110100010111)) color_data = 12'b000000001101;
		if(({row_reg, col_reg}==14'b01110100011000)) color_data = 12'b000100001011;
		if(({row_reg, col_reg}==14'b01110100011001)) color_data = 12'b001100001010;
		if(({row_reg, col_reg}==14'b01110100011010)) color_data = 12'b010000001001;
		if(({row_reg, col_reg}==14'b01110100011011)) color_data = 12'b011000001000;
		if(({row_reg, col_reg}==14'b01110100011100)) color_data = 12'b011100010111;
		if(({row_reg, col_reg}==14'b01110100011101)) color_data = 12'b100100010110;
		if(({row_reg, col_reg}==14'b01110100011110)) color_data = 12'b101100010101;
		if(({row_reg, col_reg}==14'b01110100011111)) color_data = 12'b110000100101;
		if(({row_reg, col_reg}==14'b01110100100000)) color_data = 12'b100100000010;
		if(({row_reg, col_reg}>=14'b01110100100001) && ({row_reg, col_reg}<14'b01110100100011)) color_data = 12'b100100000011;
		if(({row_reg, col_reg}==14'b01110100100011)) color_data = 12'b100000010011;
		if(({row_reg, col_reg}==14'b01110100100100)) color_data = 12'b011000010011;
		if(({row_reg, col_reg}==14'b01110100100101)) color_data = 12'b010000010010;
		if(({row_reg, col_reg}==14'b01110100100110)) color_data = 12'b010000100011;
		if(({row_reg, col_reg}==14'b01110100100111)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==14'b01110100101000)) color_data = 12'b001100010010;
		if(({row_reg, col_reg}>=14'b01110100101001) && ({row_reg, col_reg}<14'b01110100101100)) color_data = 12'b010000100011;
		if(({row_reg, col_reg}>=14'b01110100101100) && ({row_reg, col_reg}<14'b01110100110100)) color_data = 12'b010100110100;
		if(({row_reg, col_reg}==14'b01110100110100)) color_data = 12'b010100100011;
		if(({row_reg, col_reg}==14'b01110100110101)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}>=14'b01110100110110) && ({row_reg, col_reg}<14'b01110100111001)) color_data = 12'b001100010010;
		if(({row_reg, col_reg}==14'b01110100111001)) color_data = 12'b100001100111;
		if(({row_reg, col_reg}>=14'b01110100111010) && ({row_reg, col_reg}<14'b01110100111100)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==14'b01110100111100)) color_data = 12'b100101111000;
		if(({row_reg, col_reg}==14'b01110100111101)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==14'b01110100111110)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==14'b01110100111111)) color_data = 12'b101110101011;
		if(({row_reg, col_reg}==14'b01110101000000)) color_data = 12'b010000110011;
		if(({row_reg, col_reg}==14'b01110101000001)) color_data = 12'b001000000000;
		if(({row_reg, col_reg}==14'b01110101000010)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==14'b01110101000011)) color_data = 12'b110110111011;
		if(({row_reg, col_reg}==14'b01110101000100)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}>=14'b01110101000101) && ({row_reg, col_reg}<14'b01110101001010)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==14'b01110101001010)) color_data = 12'b100101111000;
		if(({row_reg, col_reg}==14'b01110101001011)) color_data = 12'b100001100111;
		if(({row_reg, col_reg}>=14'b01110101001100) && ({row_reg, col_reg}<14'b01110101001110)) color_data = 12'b010101000100;
		if(({row_reg, col_reg}>=14'b01110101001110) && ({row_reg, col_reg}<14'b01110101010001)) color_data = 12'b001100010010;
		if(({row_reg, col_reg}==14'b01110101010001)) color_data = 12'b001100010001;
		if(({row_reg, col_reg}==14'b01110101010010)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}>=14'b01110101010011) && ({row_reg, col_reg}<14'b01110101010111)) color_data = 12'b010100110100;
		if(({row_reg, col_reg}==14'b01110101010111)) color_data = 12'b001100100011;
		if(({row_reg, col_reg}==14'b01110101011000)) color_data = 12'b000000000100;
		if(({row_reg, col_reg}==14'b01110101011001)) color_data = 12'b000000001001;
		if(({row_reg, col_reg}==14'b01110101011010)) color_data = 12'b000000001101;

		if(({row_reg, col_reg}>=14'b01110101011011) && ({row_reg, col_reg}<14'b01110110010110)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==14'b01110110010110)) color_data = 12'b000000001110;
		if(({row_reg, col_reg}==14'b01110110010111)) color_data = 12'b000100001100;
		if(({row_reg, col_reg}==14'b01110110011000)) color_data = 12'b001100001001;
		if(({row_reg, col_reg}==14'b01110110011001)) color_data = 12'b011000010111;
		if(({row_reg, col_reg}==14'b01110110011010)) color_data = 12'b100000100110;
		if(({row_reg, col_reg}==14'b01110110011011)) color_data = 12'b101000100110;
		if(({row_reg, col_reg}>=14'b01110110011100) && ({row_reg, col_reg}<14'b01110110011110)) color_data = 12'b101100100101;
		if(({row_reg, col_reg}==14'b01110110011110)) color_data = 12'b110000100101;
		if(({row_reg, col_reg}==14'b01110110011111)) color_data = 12'b110000100100;
		if(({row_reg, col_reg}>=14'b01110110100000) && ({row_reg, col_reg}<14'b01110110100010)) color_data = 12'b100100000011;
		if(({row_reg, col_reg}==14'b01110110100010)) color_data = 12'b100000000011;
		if(({row_reg, col_reg}==14'b01110110100011)) color_data = 12'b100000010011;
		if(({row_reg, col_reg}==14'b01110110100100)) color_data = 12'b011000010011;
		if(({row_reg, col_reg}==14'b01110110100101)) color_data = 12'b010000010010;
		if(({row_reg, col_reg}==14'b01110110100110)) color_data = 12'b010000010011;
		if(({row_reg, col_reg}>=14'b01110110100111) && ({row_reg, col_reg}<14'b01110110101011)) color_data = 12'b001100010010;
		if(({row_reg, col_reg}==14'b01110110101011)) color_data = 12'b010000100011;
		if(({row_reg, col_reg}>=14'b01110110101100) && ({row_reg, col_reg}<14'b01110110110100)) color_data = 12'b010100110100;
		if(({row_reg, col_reg}==14'b01110110110100)) color_data = 12'b010100100011;
		if(({row_reg, col_reg}==14'b01110110110101)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}==14'b01110110110110)) color_data = 12'b001100010010;
		if(({row_reg, col_reg}==14'b01110110110111)) color_data = 12'b010000100011;
		if(({row_reg, col_reg}==14'b01110110111000)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}==14'b01110110111001)) color_data = 12'b100001100110;
		if(({row_reg, col_reg}>=14'b01110110111010) && ({row_reg, col_reg}<14'b01110110111100)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==14'b01110110111100)) color_data = 12'b100101111000;
		if(({row_reg, col_reg}==14'b01110110111101)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==14'b01110110111110)) color_data = 12'b110010101011;
		if(({row_reg, col_reg}==14'b01110110111111)) color_data = 12'b110010111011;
		if(({row_reg, col_reg}==14'b01110111000000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==14'b01110111000001)) color_data = 12'b001000000000;
		if(({row_reg, col_reg}==14'b01110111000010)) color_data = 12'b100001100110;
		if(({row_reg, col_reg}==14'b01110111000011)) color_data = 12'b110110111011;
		if(({row_reg, col_reg}==14'b01110111000100)) color_data = 12'b101110011001;
		if(({row_reg, col_reg}>=14'b01110111000101) && ({row_reg, col_reg}<14'b01110111001001)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==14'b01110111001001)) color_data = 12'b100101111000;
		if(({row_reg, col_reg}==14'b01110111001010)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==14'b01110111001011)) color_data = 12'b100001100111;
		if(({row_reg, col_reg}==14'b01110111001100)) color_data = 12'b010000100011;
		if(({row_reg, col_reg}==14'b01110111001101)) color_data = 12'b010100110100;
		if(({row_reg, col_reg}==14'b01110111001110)) color_data = 12'b001100010010;
		if(({row_reg, col_reg}==14'b01110111001111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=14'b01110111010000) && ({row_reg, col_reg}<14'b01110111010010)) color_data = 12'b001100010010;
		if(({row_reg, col_reg}==14'b01110111010010)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}>=14'b01110111010011) && ({row_reg, col_reg}<14'b01110111010111)) color_data = 12'b010100110100;
		if(({row_reg, col_reg}==14'b01110111010111)) color_data = 12'b001100100100;
		if(({row_reg, col_reg}==14'b01110111011000)) color_data = 12'b000000000101;
		if(({row_reg, col_reg}==14'b01110111011001)) color_data = 12'b000000001001;
		if(({row_reg, col_reg}==14'b01110111011010)) color_data = 12'b000000001101;

		if(({row_reg, col_reg}>=14'b01110111011011) && ({row_reg, col_reg}<14'b01111000010110)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==14'b01111000010110)) color_data = 12'b000100001101;
		if(({row_reg, col_reg}==14'b01111000010111)) color_data = 12'b001000001011;
		if(({row_reg, col_reg}==14'b01111000011000)) color_data = 12'b010100001000;
		if(({row_reg, col_reg}==14'b01111000011001)) color_data = 12'b100000010111;
		if(({row_reg, col_reg}==14'b01111000011010)) color_data = 12'b101000100101;
		if(({row_reg, col_reg}>=14'b01111000011011) && ({row_reg, col_reg}<14'b01111000011101)) color_data = 12'b101000010100;
		if(({row_reg, col_reg}==14'b01111000011101)) color_data = 12'b100100010011;
		if(({row_reg, col_reg}>=14'b01111000011110) && ({row_reg, col_reg}<14'b01111000100001)) color_data = 12'b100100010100;
		if(({row_reg, col_reg}==14'b01111000100001)) color_data = 12'b100100000100;
		if(({row_reg, col_reg}==14'b01111000100010)) color_data = 12'b100000000011;
		if(({row_reg, col_reg}==14'b01111000100011)) color_data = 12'b100000010011;
		if(({row_reg, col_reg}==14'b01111000100100)) color_data = 12'b011000010010;
		if(({row_reg, col_reg}==14'b01111000100101)) color_data = 12'b010100010010;
		if(({row_reg, col_reg}>=14'b01111000100110) && ({row_reg, col_reg}<14'b01111000101000)) color_data = 12'b010000010010;
		if(({row_reg, col_reg}>=14'b01111000101000) && ({row_reg, col_reg}<14'b01111000101011)) color_data = 12'b001100010010;
		if(({row_reg, col_reg}>=14'b01111000101011) && ({row_reg, col_reg}<14'b01111000101110)) color_data = 12'b010000100011;
		if(({row_reg, col_reg}>=14'b01111000101110) && ({row_reg, col_reg}<14'b01111000110000)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}>=14'b01111000110000) && ({row_reg, col_reg}<14'b01111000110100)) color_data = 12'b010000100011;
		if(({row_reg, col_reg}>=14'b01111000110100) && ({row_reg, col_reg}<14'b01111000110111)) color_data = 12'b001100010010;
		if(({row_reg, col_reg}==14'b01111000110111)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}==14'b01111000111000)) color_data = 12'b001100010010;
		if(({row_reg, col_reg}==14'b01111000111001)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==14'b01111000111010)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}>=14'b01111000111011) && ({row_reg, col_reg}<14'b01111000111101)) color_data = 12'b100101111000;
		if(({row_reg, col_reg}>=14'b01111000111101) && ({row_reg, col_reg}<14'b01111001000000)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==14'b01111001000000)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}==14'b01111001000001)) color_data = 12'b001000000000;
		if(({row_reg, col_reg}==14'b01111001000010)) color_data = 12'b100001100110;
		if(({row_reg, col_reg}==14'b01111001000011)) color_data = 12'b110110111011;
		if(({row_reg, col_reg}==14'b01111001000100)) color_data = 12'b101110011001;
		if(({row_reg, col_reg}>=14'b01111001000101) && ({row_reg, col_reg}<14'b01111001001000)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==14'b01111001001000)) color_data = 12'b100101111000;
		if(({row_reg, col_reg}==14'b01111001001001)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==14'b01111001001010)) color_data = 12'b101010001001;
		if(({row_reg, col_reg}==14'b01111001001011)) color_data = 12'b100001100111;
		if(({row_reg, col_reg}==14'b01111001001100)) color_data = 12'b001100010010;
		if(({row_reg, col_reg}==14'b01111001001101)) color_data = 12'b010000100011;
		if(({row_reg, col_reg}>=14'b01111001001110) && ({row_reg, col_reg}<14'b01111001010000)) color_data = 12'b001100010010;
		if(({row_reg, col_reg}>=14'b01111001010000) && ({row_reg, col_reg}<14'b01111001010010)) color_data = 12'b001100010001;
		if(({row_reg, col_reg}==14'b01111001010010)) color_data = 12'b001100010010;
		if(({row_reg, col_reg}>=14'b01111001010011) && ({row_reg, col_reg}<14'b01111001010101)) color_data = 12'b010000100011;
		if(({row_reg, col_reg}>=14'b01111001010101) && ({row_reg, col_reg}<14'b01111001010111)) color_data = 12'b001100010010;
		if(({row_reg, col_reg}==14'b01111001010111)) color_data = 12'b001100010011;
		if(({row_reg, col_reg}==14'b01111001011000)) color_data = 12'b000000000101;
		if(({row_reg, col_reg}==14'b01111001011001)) color_data = 12'b000000001010;
		if(({row_reg, col_reg}==14'b01111001011010)) color_data = 12'b000000001110;

		if(({row_reg, col_reg}>=14'b01111001011011) && ({row_reg, col_reg}<14'b01111010010110)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==14'b01111010010110)) color_data = 12'b000100001101;
		if(({row_reg, col_reg}==14'b01111010010111)) color_data = 12'b001000001011;
		if(({row_reg, col_reg}==14'b01111010011000)) color_data = 12'b010000001001;
		if(({row_reg, col_reg}==14'b01111010011001)) color_data = 12'b011000000111;
		if(({row_reg, col_reg}==14'b01111010011010)) color_data = 12'b011100010110;
		if(({row_reg, col_reg}==14'b01111010011011)) color_data = 12'b011100000101;
		if(({row_reg, col_reg}>=14'b01111010011100) && ({row_reg, col_reg}<14'b01111010100000)) color_data = 12'b011000000101;
		if(({row_reg, col_reg}>=14'b01111010100000) && ({row_reg, col_reg}<14'b01111010100010)) color_data = 12'b100000000100;
		if(({row_reg, col_reg}>=14'b01111010100010) && ({row_reg, col_reg}<14'b01111010100100)) color_data = 12'b100000010011;
		if(({row_reg, col_reg}==14'b01111010100100)) color_data = 12'b011000010010;
		if(({row_reg, col_reg}==14'b01111010100101)) color_data = 12'b010100000010;
		if(({row_reg, col_reg}==14'b01111010100110)) color_data = 12'b010000010010;
		if(({row_reg, col_reg}==14'b01111010100111)) color_data = 12'b010000010011;
		if(({row_reg, col_reg}>=14'b01111010101000) && ({row_reg, col_reg}<14'b01111010101100)) color_data = 12'b001100010010;
		if(({row_reg, col_reg}==14'b01111010101100)) color_data = 12'b010000010010;
		if(({row_reg, col_reg}>=14'b01111010101101) && ({row_reg, col_reg}<14'b01111010110000)) color_data = 12'b001100010010;
		if(({row_reg, col_reg}==14'b01111010110000)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}>=14'b01111010110001) && ({row_reg, col_reg}<14'b01111010110011)) color_data = 12'b001100010010;
		if(({row_reg, col_reg}==14'b01111010110011)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}>=14'b01111010110100) && ({row_reg, col_reg}<14'b01111010110111)) color_data = 12'b001100010010;
		if(({row_reg, col_reg}==14'b01111010110111)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==14'b01111010111000)) color_data = 12'b001100010001;
		if(({row_reg, col_reg}==14'b01111010111001)) color_data = 12'b100001100111;
		if(({row_reg, col_reg}==14'b01111010111010)) color_data = 12'b101010001001;
		if(({row_reg, col_reg}==14'b01111010111011)) color_data = 12'b100101111000;
		if(({row_reg, col_reg}>=14'b01111010111100) && ({row_reg, col_reg}<14'b01111011000000)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==14'b01111011000000)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}==14'b01111011000001)) color_data = 12'b001000000000;
		if(({row_reg, col_reg}==14'b01111011000010)) color_data = 12'b100001100110;
		if(({row_reg, col_reg}==14'b01111011000011)) color_data = 12'b110110111011;
		if(({row_reg, col_reg}==14'b01111011000100)) color_data = 12'b101110011001;
		if(({row_reg, col_reg}>=14'b01111011000101) && ({row_reg, col_reg}<14'b01111011001001)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==14'b01111011001001)) color_data = 12'b100110001001;
		if(({row_reg, col_reg}==14'b01111011001010)) color_data = 12'b101010001001;
		if(({row_reg, col_reg}==14'b01111011001011)) color_data = 12'b011101010110;
		if(({row_reg, col_reg}==14'b01111011001100)) color_data = 12'b001000000001;
		if(({row_reg, col_reg}==14'b01111011001101)) color_data = 12'b001100010010;
		if(({row_reg, col_reg}==14'b01111011001110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=14'b01111011001111) && ({row_reg, col_reg}<14'b01111011010010)) color_data = 12'b001100010010;
		if(({row_reg, col_reg}==14'b01111011010010)) color_data = 12'b001100010001;
		if(({row_reg, col_reg}>=14'b01111011010011) && ({row_reg, col_reg}<14'b01111011010111)) color_data = 12'b001100010010;
		if(({row_reg, col_reg}==14'b01111011010111)) color_data = 12'b001100100100;
		if(({row_reg, col_reg}==14'b01111011011000)) color_data = 12'b000000000101;
		if(({row_reg, col_reg}==14'b01111011011001)) color_data = 12'b000000001010;
		if(({row_reg, col_reg}==14'b01111011011010)) color_data = 12'b000000001110;

		if(({row_reg, col_reg}>=14'b01111011011011) && ({row_reg, col_reg}<14'b01111100010110)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==14'b01111100010110)) color_data = 12'b000000001110;
		if(({row_reg, col_reg}==14'b01111100010111)) color_data = 12'b000100001100;
		if(({row_reg, col_reg}==14'b01111100011000)) color_data = 12'b001000001011;
		if(({row_reg, col_reg}==14'b01111100011001)) color_data = 12'b001100001010;
		if(({row_reg, col_reg}==14'b01111100011010)) color_data = 12'b010000001010;
		if(({row_reg, col_reg}>=14'b01111100011011) && ({row_reg, col_reg}<14'b01111100011101)) color_data = 12'b001100001010;
		if(({row_reg, col_reg}>=14'b01111100011101) && ({row_reg, col_reg}<14'b01111100011111)) color_data = 12'b001100001001;
		if(({row_reg, col_reg}==14'b01111100011111)) color_data = 12'b010000001000;
		if(({row_reg, col_reg}==14'b01111100100000)) color_data = 12'b011100000100;
		if(({row_reg, col_reg}==14'b01111100100001)) color_data = 12'b100000000100;
		if(({row_reg, col_reg}==14'b01111100100010)) color_data = 12'b100000010100;
		if(({row_reg, col_reg}==14'b01111100100011)) color_data = 12'b100000010011;
		if(({row_reg, col_reg}==14'b01111100100100)) color_data = 12'b011100010011;
		if(({row_reg, col_reg}==14'b01111100100101)) color_data = 12'b011000010011;
		if(({row_reg, col_reg}==14'b01111100100110)) color_data = 12'b010100010011;
		if(({row_reg, col_reg}==14'b01111100100111)) color_data = 12'b010000010011;
		if(({row_reg, col_reg}==14'b01111100101000)) color_data = 12'b001100010010;
		if(({row_reg, col_reg}>=14'b01111100101001) && ({row_reg, col_reg}<14'b01111100101011)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}>=14'b01111100101011) && ({row_reg, col_reg}<14'b01111100101101)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}==14'b01111100101101)) color_data = 12'b010000010010;
		if(({row_reg, col_reg}==14'b01111100101110)) color_data = 12'b010000100011;
		if(({row_reg, col_reg}==14'b01111100101111)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}>=14'b01111100110000) && ({row_reg, col_reg}<14'b01111100110011)) color_data = 12'b001100010010;
		if(({row_reg, col_reg}==14'b01111100110011)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==14'b01111100110100)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}>=14'b01111100110101) && ({row_reg, col_reg}<14'b01111100110111)) color_data = 12'b001100010010;
		if(({row_reg, col_reg}==14'b01111100110111)) color_data = 12'b010100110100;
		if(({row_reg, col_reg}==14'b01111100111000)) color_data = 12'b010100110011;
		if(({row_reg, col_reg}==14'b01111100111001)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==14'b01111100111010)) color_data = 12'b101010001000;
		if(({row_reg, col_reg}>=14'b01111100111011) && ({row_reg, col_reg}<14'b01111100111110)) color_data = 12'b100101111000;
		if(({row_reg, col_reg}>=14'b01111100111110) && ({row_reg, col_reg}<14'b01111101000000)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==14'b01111101000000)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}==14'b01111101000001)) color_data = 12'b001000000000;
		if(({row_reg, col_reg}==14'b01111101000010)) color_data = 12'b100001100110;
		if(({row_reg, col_reg}==14'b01111101000011)) color_data = 12'b110110111011;
		if(({row_reg, col_reg}==14'b01111101000100)) color_data = 12'b101110011010;
		if(({row_reg, col_reg}>=14'b01111101000101) && ({row_reg, col_reg}<14'b01111101000111)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}>=14'b01111101000111) && ({row_reg, col_reg}<14'b01111101001001)) color_data = 12'b100101111000;
		if(({row_reg, col_reg}==14'b01111101001001)) color_data = 12'b100001111000;
		if(({row_reg, col_reg}==14'b01111101001010)) color_data = 12'b100001100111;
		if(({row_reg, col_reg}==14'b01111101001011)) color_data = 12'b011101010110;
		if(({row_reg, col_reg}==14'b01111101001100)) color_data = 12'b010000100011;
		if(({row_reg, col_reg}==14'b01111101001101)) color_data = 12'b010100110011;
		if(({row_reg, col_reg}>=14'b01111101001110) && ({row_reg, col_reg}<14'b01111101010010)) color_data = 12'b001100010010;
		if(({row_reg, col_reg}==14'b01111101010010)) color_data = 12'b001100010001;
		if(({row_reg, col_reg}>=14'b01111101010011) && ({row_reg, col_reg}<14'b01111101010111)) color_data = 12'b001100010010;
		if(({row_reg, col_reg}==14'b01111101010111)) color_data = 12'b001000010011;
		if(({row_reg, col_reg}==14'b01111101011000)) color_data = 12'b000000000101;
		if(({row_reg, col_reg}==14'b01111101011001)) color_data = 12'b000000001010;
		if(({row_reg, col_reg}==14'b01111101011010)) color_data = 12'b000000001110;

		if(({row_reg, col_reg}>=14'b01111101011011) && ({row_reg, col_reg}<14'b01111110010111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==14'b01111110010111)) color_data = 12'b000000001110;
		if(({row_reg, col_reg}>=14'b01111110011000) && ({row_reg, col_reg}<14'b01111110011011)) color_data = 12'b000100001101;
		if(({row_reg, col_reg}==14'b01111110011011)) color_data = 12'b000000001101;
		if(({row_reg, col_reg}>=14'b01111110011100) && ({row_reg, col_reg}<14'b01111110011110)) color_data = 12'b000100001101;
		if(({row_reg, col_reg}==14'b01111110011110)) color_data = 12'b001000001011;
		if(({row_reg, col_reg}==14'b01111110011111)) color_data = 12'b001000001010;
		if(({row_reg, col_reg}>=14'b01111110100000) && ({row_reg, col_reg}<14'b01111110100010)) color_data = 12'b011100000100;
		if(({row_reg, col_reg}==14'b01111110100010)) color_data = 12'b100000000100;
		if(({row_reg, col_reg}==14'b01111110100011)) color_data = 12'b100000000011;
		if(({row_reg, col_reg}==14'b01111110100100)) color_data = 12'b011100010011;
		if(({row_reg, col_reg}==14'b01111110100101)) color_data = 12'b011100010100;
		if(({row_reg, col_reg}==14'b01111110100110)) color_data = 12'b011000010011;
		if(({row_reg, col_reg}==14'b01111110100111)) color_data = 12'b010000010011;
		if(({row_reg, col_reg}==14'b01111110101000)) color_data = 12'b001100010010;
		if(({row_reg, col_reg}>=14'b01111110101001) && ({row_reg, col_reg}<14'b01111110101100)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==14'b01111110101100)) color_data = 12'b010000010010;
		if(({row_reg, col_reg}==14'b01111110101101)) color_data = 12'b001100010010;
		if(({row_reg, col_reg}>=14'b01111110101110) && ({row_reg, col_reg}<14'b01111110110000)) color_data = 12'b001100010011;
		if(({row_reg, col_reg}==14'b01111110110000)) color_data = 12'b001100010010;
		if(({row_reg, col_reg}>=14'b01111110110001) && ({row_reg, col_reg}<14'b01111110110011)) color_data = 12'b001100100011;
		if(({row_reg, col_reg}>=14'b01111110110011) && ({row_reg, col_reg}<14'b01111110110110)) color_data = 12'b001100010010;
		if(({row_reg, col_reg}==14'b01111110110110)) color_data = 12'b010000100011;
		if(({row_reg, col_reg}==14'b01111110110111)) color_data = 12'b100001100110;
		if(({row_reg, col_reg}==14'b01111110111000)) color_data = 12'b011101010110;
		if(({row_reg, col_reg}==14'b01111110111001)) color_data = 12'b100101110111;
		if(({row_reg, col_reg}>=14'b01111110111010) && ({row_reg, col_reg}<14'b01111110111100)) color_data = 12'b100101111000;
		if(({row_reg, col_reg}==14'b01111110111100)) color_data = 12'b101010001000;
		if(({row_reg, col_reg}>=14'b01111110111101) && ({row_reg, col_reg}<14'b01111111000000)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==14'b01111111000000)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}==14'b01111111000001)) color_data = 12'b001000000000;
		if(({row_reg, col_reg}==14'b01111111000010)) color_data = 12'b100001100110;
		if(({row_reg, col_reg}==14'b01111111000011)) color_data = 12'b110110111011;
		if(({row_reg, col_reg}==14'b01111111000100)) color_data = 12'b101110011010;
		if(({row_reg, col_reg}>=14'b01111111000101) && ({row_reg, col_reg}<14'b01111111000111)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}>=14'b01111111000111) && ({row_reg, col_reg}<14'b01111111001001)) color_data = 12'b100101111000;
		if(({row_reg, col_reg}==14'b01111111001001)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==14'b01111111001010)) color_data = 12'b011001010101;
		if(({row_reg, col_reg}>=14'b01111111001011) && ({row_reg, col_reg}<14'b01111111001110)) color_data = 12'b011101010110;
		if(({row_reg, col_reg}==14'b01111111001110)) color_data = 12'b001100010010;
		if(({row_reg, col_reg}==14'b01111111001111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==14'b01111111010000)) color_data = 12'b001100010010;
		if(({row_reg, col_reg}>=14'b01111111010001) && ({row_reg, col_reg}<14'b01111111010011)) color_data = 12'b001100010001;
		if(({row_reg, col_reg}>=14'b01111111010011) && ({row_reg, col_reg}<14'b01111111010111)) color_data = 12'b001100010010;
		if(({row_reg, col_reg}==14'b01111111010111)) color_data = 12'b001000010010;
		if(({row_reg, col_reg}==14'b01111111011000)) color_data = 12'b000000000101;
		if(({row_reg, col_reg}==14'b01111111011001)) color_data = 12'b000000001001;
		if(({row_reg, col_reg}==14'b01111111011010)) color_data = 12'b000000001110;

		if(({row_reg, col_reg}>=14'b01111111011011) && ({row_reg, col_reg}<14'b10000000011101)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==14'b10000000011101)) color_data = 12'b000000001110;
		if(({row_reg, col_reg}==14'b10000000011110)) color_data = 12'b000100001101;
		if(({row_reg, col_reg}==14'b10000000011111)) color_data = 12'b001000001100;
		if(({row_reg, col_reg}==14'b10000000100000)) color_data = 12'b011000000101;
		if(({row_reg, col_reg}==14'b10000000100001)) color_data = 12'b100000010101;
		if(({row_reg, col_reg}==14'b10000000100010)) color_data = 12'b100100000011;
		if(({row_reg, col_reg}==14'b10000000100011)) color_data = 12'b100100010010;
		if(({row_reg, col_reg}==14'b10000000100100)) color_data = 12'b100100010011;
		if(({row_reg, col_reg}==14'b10000000100101)) color_data = 12'b011100010100;
		if(({row_reg, col_reg}==14'b10000000100110)) color_data = 12'b010100010110;
		if(({row_reg, col_reg}==14'b10000000100111)) color_data = 12'b001100000110;
		if(({row_reg, col_reg}==14'b10000000101000)) color_data = 12'b001100000101;
		if(({row_reg, col_reg}==14'b10000000101001)) color_data = 12'b001100000100;
		if(({row_reg, col_reg}==14'b10000000101010)) color_data = 12'b001100010011;
		if(({row_reg, col_reg}>=14'b10000000101011) && ({row_reg, col_reg}<14'b10000000101101)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==14'b10000000101101)) color_data = 12'b001100010010;
		if(({row_reg, col_reg}>=14'b10000000101110) && ({row_reg, col_reg}<14'b10000000110000)) color_data = 12'b001100010011;
		if(({row_reg, col_reg}==14'b10000000110000)) color_data = 12'b001100010001;
		if(({row_reg, col_reg}==14'b10000000110001)) color_data = 12'b001100010010;
		if(({row_reg, col_reg}==14'b10000000110010)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}==14'b10000000110011)) color_data = 12'b001100010010;
		if(({row_reg, col_reg}>=14'b10000000110100) && ({row_reg, col_reg}<14'b10000000110110)) color_data = 12'b010000100011;
		if(({row_reg, col_reg}==14'b10000000110110)) color_data = 12'b010000110011;
		if(({row_reg, col_reg}>=14'b10000000110111) && ({row_reg, col_reg}<14'b10000000111001)) color_data = 12'b011101010101;
		if(({row_reg, col_reg}==14'b10000000111001)) color_data = 12'b100001100111;
		if(({row_reg, col_reg}==14'b10000000111010)) color_data = 12'b101010001000;
		if(({row_reg, col_reg}==14'b10000000111011)) color_data = 12'b100101111000;
		if(({row_reg, col_reg}==14'b10000000111100)) color_data = 12'b100001100110;
		if(({row_reg, col_reg}==14'b10000000111101)) color_data = 12'b100101110111;
		if(({row_reg, col_reg}==14'b10000000111110)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==14'b10000000111111)) color_data = 12'b100001100110;
		if(({row_reg, col_reg}==14'b10000001000000)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==14'b10000001000001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==14'b10000001000010)) color_data = 12'b011101010110;
		if(({row_reg, col_reg}==14'b10000001000011)) color_data = 12'b101110011010;
		if(({row_reg, col_reg}>=14'b10000001000100) && ({row_reg, col_reg}<14'b10000001000110)) color_data = 12'b101010001000;
		if(({row_reg, col_reg}==14'b10000001000110)) color_data = 12'b100101111000;
		if(({row_reg, col_reg}>=14'b10000001000111) && ({row_reg, col_reg}<14'b10000001001001)) color_data = 12'b100101111001;
		if(({row_reg, col_reg}==14'b10000001001001)) color_data = 12'b100001100111;
		if(({row_reg, col_reg}==14'b10000001001010)) color_data = 12'b011101010110;
		if(({row_reg, col_reg}>=14'b10000001001011) && ({row_reg, col_reg}<14'b10000001001101)) color_data = 12'b011101010101;
		if(({row_reg, col_reg}==14'b10000001001101)) color_data = 12'b011001000100;
		if(({row_reg, col_reg}==14'b10000001001110)) color_data = 12'b010000100011;
		if(({row_reg, col_reg}==14'b10000001001111)) color_data = 12'b010000010011;
		if(({row_reg, col_reg}>=14'b10000001010000) && ({row_reg, col_reg}<14'b10000001010100)) color_data = 12'b001100010001;
		if(({row_reg, col_reg}==14'b10000001010100)) color_data = 12'b001100010010;
		if(({row_reg, col_reg}==14'b10000001010101)) color_data = 12'b001000010011;
		if(({row_reg, col_reg}==14'b10000001010110)) color_data = 12'b000100000100;
		if(({row_reg, col_reg}==14'b10000001010111)) color_data = 12'b000000000111;
		if(({row_reg, col_reg}==14'b10000001011000)) color_data = 12'b000000001010;
		if(({row_reg, col_reg}==14'b10000001011001)) color_data = 12'b000000001101;
		if(({row_reg, col_reg}==14'b10000001011010)) color_data = 12'b000000001110;

		if(({row_reg, col_reg}>=14'b10000001011011) && ({row_reg, col_reg}<14'b10000010011101)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==14'b10000010011101)) color_data = 12'b000000001110;
		if(({row_reg, col_reg}==14'b10000010011110)) color_data = 12'b000100001100;
		if(({row_reg, col_reg}==14'b10000010011111)) color_data = 12'b001000001011;
		if(({row_reg, col_reg}==14'b10000010100000)) color_data = 12'b011100000100;
		if(({row_reg, col_reg}==14'b10000010100001)) color_data = 12'b101000100101;
		if(({row_reg, col_reg}==14'b10000010100010)) color_data = 12'b101100100100;
		if(({row_reg, col_reg}==14'b10000010100011)) color_data = 12'b101000100100;
		if(({row_reg, col_reg}==14'b10000010100100)) color_data = 12'b100100010101;
		if(({row_reg, col_reg}==14'b10000010100101)) color_data = 12'b011000000101;
		if(({row_reg, col_reg}==14'b10000010100110)) color_data = 12'b010000000111;
		if(({row_reg, col_reg}==14'b10000010100111)) color_data = 12'b001000001000;
		if(({row_reg, col_reg}==14'b10000010101000)) color_data = 12'b001000000111;
		if(({row_reg, col_reg}==14'b10000010101001)) color_data = 12'b001000000110;
		if(({row_reg, col_reg}==14'b10000010101010)) color_data = 12'b001000000100;
		if(({row_reg, col_reg}==14'b10000010101011)) color_data = 12'b001000010011;
		if(({row_reg, col_reg}>=14'b10000010101100) && ({row_reg, col_reg}<14'b10000010110000)) color_data = 12'b001100010010;
		if(({row_reg, col_reg}==14'b10000010110000)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}>=14'b10000010110001) && ({row_reg, col_reg}<14'b10000010110100)) color_data = 12'b001100010010;
		if(({row_reg, col_reg}==14'b10000010110100)) color_data = 12'b010100110100;
		if(({row_reg, col_reg}>=14'b10000010110101) && ({row_reg, col_reg}<14'b10000010110111)) color_data = 12'b011101010110;
		if(({row_reg, col_reg}==14'b10000010110111)) color_data = 12'b100001100110;
		if(({row_reg, col_reg}==14'b10000010111000)) color_data = 12'b011101010110;
		if(({row_reg, col_reg}==14'b10000010111001)) color_data = 12'b100101110111;
		if(({row_reg, col_reg}==14'b10000010111010)) color_data = 12'b100101111000;
		if(({row_reg, col_reg}==14'b10000010111011)) color_data = 12'b011001000101;
		if(({row_reg, col_reg}==14'b10000010111100)) color_data = 12'b001000000001;
		if(({row_reg, col_reg}>=14'b10000010111101) && ({row_reg, col_reg}<14'b10000011000001)) color_data = 12'b001100010001;
		if(({row_reg, col_reg}==14'b10000011000001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=14'b10000011000010) && ({row_reg, col_reg}<14'b10000011000100)) color_data = 12'b001100010001;
		if(({row_reg, col_reg}==14'b10000011000100)) color_data = 12'b010000110011;
		if(({row_reg, col_reg}==14'b10000011000101)) color_data = 12'b100101110111;
		if(({row_reg, col_reg}>=14'b10000011000110) && ({row_reg, col_reg}<14'b10000011001000)) color_data = 12'b100101111000;
		if(({row_reg, col_reg}==14'b10000011001000)) color_data = 12'b100101111001;
		if(({row_reg, col_reg}==14'b10000011001001)) color_data = 12'b100001100111;
		if(({row_reg, col_reg}>=14'b10000011001010) && ({row_reg, col_reg}<14'b10000011001100)) color_data = 12'b011101010110;
		if(({row_reg, col_reg}>=14'b10000011001100) && ({row_reg, col_reg}<14'b10000011001110)) color_data = 12'b011101010101;
		if(({row_reg, col_reg}==14'b10000011001110)) color_data = 12'b011101010110;
		if(({row_reg, col_reg}==14'b10000011001111)) color_data = 12'b011101010111;
		if(({row_reg, col_reg}==14'b10000011010000)) color_data = 12'b001100100011;
		if(({row_reg, col_reg}==14'b10000011010001)) color_data = 12'b001100010011;
		if(({row_reg, col_reg}>=14'b10000011010010) && ({row_reg, col_reg}<14'b10000011010100)) color_data = 12'b001100010100;
		if(({row_reg, col_reg}==14'b10000011010100)) color_data = 12'b001000010100;
		if(({row_reg, col_reg}==14'b10000011010101)) color_data = 12'b000100000100;
		if(({row_reg, col_reg}==14'b10000011010110)) color_data = 12'b000000000110;
		if(({row_reg, col_reg}==14'b10000011010111)) color_data = 12'b000000001001;
		if(({row_reg, col_reg}==14'b10000011011000)) color_data = 12'b000000001011;
		if(({row_reg, col_reg}==14'b10000011011001)) color_data = 12'b000000001101;

		if(({row_reg, col_reg}>=14'b10000011011010) && ({row_reg, col_reg}<14'b10000100011101)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==14'b10000100011101)) color_data = 12'b000100001101;
		if(({row_reg, col_reg}==14'b10000100011110)) color_data = 12'b001000001011;
		if(({row_reg, col_reg}==14'b10000100011111)) color_data = 12'b001100001011;
		if(({row_reg, col_reg}==14'b10000100100000)) color_data = 12'b100100010100;
		if(({row_reg, col_reg}==14'b10000100100001)) color_data = 12'b101100110110;
		if(({row_reg, col_reg}==14'b10000100100010)) color_data = 12'b101100110101;
		if(({row_reg, col_reg}==14'b10000100100011)) color_data = 12'b101000100101;
		if(({row_reg, col_reg}==14'b10000100100100)) color_data = 12'b100000010110;
		if(({row_reg, col_reg}==14'b10000100100101)) color_data = 12'b010000001000;
		if(({row_reg, col_reg}==14'b10000100100110)) color_data = 12'b001000001001;
		if(({row_reg, col_reg}==14'b10000100100111)) color_data = 12'b000100001011;
		if(({row_reg, col_reg}==14'b10000100101000)) color_data = 12'b000000001010;
		if(({row_reg, col_reg}==14'b10000100101001)) color_data = 12'b000000001001;
		if(({row_reg, col_reg}==14'b10000100101010)) color_data = 12'b000100000110;
		if(({row_reg, col_reg}==14'b10000100101011)) color_data = 12'b000100000100;
		if(({row_reg, col_reg}==14'b10000100101100)) color_data = 12'b001000010011;
		if(({row_reg, col_reg}==14'b10000100101101)) color_data = 12'b001100010011;
		if(({row_reg, col_reg}>=14'b10000100101110) && ({row_reg, col_reg}<14'b10000100110000)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}>=14'b10000100110000) && ({row_reg, col_reg}<14'b10000100110100)) color_data = 12'b001100010010;
		if(({row_reg, col_reg}==14'b10000100110100)) color_data = 12'b010100110100;
		if(({row_reg, col_reg}>=14'b10000100110101) && ({row_reg, col_reg}<14'b10000100111001)) color_data = 12'b011101010110;
		if(({row_reg, col_reg}==14'b10000100111001)) color_data = 12'b100101111000;
		if(({row_reg, col_reg}==14'b10000100111010)) color_data = 12'b101001111001;
		if(({row_reg, col_reg}==14'b10000100111011)) color_data = 12'b011001000101;
		if(({row_reg, col_reg}==14'b10000100111100)) color_data = 12'b001100010001;
		if(({row_reg, col_reg}==14'b10000100111101)) color_data = 12'b001100010010;
		if(({row_reg, col_reg}==14'b10000100111110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==14'b10000100111111)) color_data = 12'b001100010001;
		if(({row_reg, col_reg}==14'b10000101000000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==14'b10000101000001)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==14'b10000101000010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==14'b10000101000011)) color_data = 12'b001000000000;
		if(({row_reg, col_reg}==14'b10000101000100)) color_data = 12'b010100110011;
		if(({row_reg, col_reg}==14'b10000101000101)) color_data = 12'b101010001000;
		if(({row_reg, col_reg}>=14'b10000101000110) && ({row_reg, col_reg}<14'b10000101001000)) color_data = 12'b100101111000;
		if(({row_reg, col_reg}==14'b10000101001000)) color_data = 12'b100101111001;
		if(({row_reg, col_reg}==14'b10000101001001)) color_data = 12'b100001101000;
		if(({row_reg, col_reg}==14'b10000101001010)) color_data = 12'b011101010111;
		if(({row_reg, col_reg}>=14'b10000101001011) && ({row_reg, col_reg}<14'b10000101001110)) color_data = 12'b011101010110;
		if(({row_reg, col_reg}>=14'b10000101001110) && ({row_reg, col_reg}<14'b10000101010000)) color_data = 12'b011101010111;
		if(({row_reg, col_reg}==14'b10000101010000)) color_data = 12'b000100010101;
		if(({row_reg, col_reg}>=14'b10000101010001) && ({row_reg, col_reg}<14'b10000101010011)) color_data = 12'b000000000101;
		if(({row_reg, col_reg}>=14'b10000101010011) && ({row_reg, col_reg}<14'b10000101010101)) color_data = 12'b000000000110;
		if(({row_reg, col_reg}==14'b10000101010101)) color_data = 12'b000000000111;
		if(({row_reg, col_reg}==14'b10000101010110)) color_data = 12'b000000001000;
		if(({row_reg, col_reg}==14'b10000101010111)) color_data = 12'b000000001011;
		if(({row_reg, col_reg}==14'b10000101011000)) color_data = 12'b000000001101;
		if(({row_reg, col_reg}==14'b10000101011001)) color_data = 12'b000000001110;

		if(({row_reg, col_reg}>=14'b10000101011010) && ({row_reg, col_reg}<14'b10000110011100)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==14'b10000110011100)) color_data = 12'b000000001110;
		if(({row_reg, col_reg}==14'b10000110011101)) color_data = 12'b000100001100;
		if(({row_reg, col_reg}==14'b10000110011110)) color_data = 12'b001100001011;
		if(({row_reg, col_reg}==14'b10000110011111)) color_data = 12'b010000001010;
		if(({row_reg, col_reg}==14'b10000110100000)) color_data = 12'b100100010101;
		if(({row_reg, col_reg}==14'b10000110100001)) color_data = 12'b101000100110;
		if(({row_reg, col_reg}==14'b10000110100010)) color_data = 12'b100100010101;
		if(({row_reg, col_reg}==14'b10000110100011)) color_data = 12'b011100000110;
		if(({row_reg, col_reg}==14'b10000110100100)) color_data = 12'b010100001000;
		if(({row_reg, col_reg}==14'b10000110100101)) color_data = 12'b001100001010;
		if(({row_reg, col_reg}==14'b10000110100110)) color_data = 12'b000100001100;
		if(({row_reg, col_reg}>=14'b10000110100111) && ({row_reg, col_reg}<14'b10000110101001)) color_data = 12'b000000001110;
		if(({row_reg, col_reg}==14'b10000110101001)) color_data = 12'b000000001100;
		if(({row_reg, col_reg}==14'b10000110101010)) color_data = 12'b000000001001;
		if(({row_reg, col_reg}==14'b10000110101011)) color_data = 12'b000000000111;
		if(({row_reg, col_reg}==14'b10000110101100)) color_data = 12'b000100000101;
		if(({row_reg, col_reg}==14'b10000110101101)) color_data = 12'b001000010100;
		if(({row_reg, col_reg}==14'b10000110101110)) color_data = 12'b001100010011;
		if(({row_reg, col_reg}==14'b10000110101111)) color_data = 12'b001100010010;
		if(({row_reg, col_reg}>=14'b10000110110000) && ({row_reg, col_reg}<14'b10000110110010)) color_data = 12'b001100010011;
		if(({row_reg, col_reg}==14'b10000110110010)) color_data = 12'b010101000100;
		if(({row_reg, col_reg}==14'b10000110110011)) color_data = 12'b011101000101;
		if(({row_reg, col_reg}==14'b10000110110100)) color_data = 12'b011101010101;
		if(({row_reg, col_reg}==14'b10000110110101)) color_data = 12'b100001010110;
		if(({row_reg, col_reg}==14'b10000110110110)) color_data = 12'b011101010111;
		if(({row_reg, col_reg}==14'b10000110110111)) color_data = 12'b100001010111;
		if(({row_reg, col_reg}==14'b10000110111000)) color_data = 12'b011101010111;
		if(({row_reg, col_reg}==14'b10000110111001)) color_data = 12'b100101101000;
		if(({row_reg, col_reg}==14'b10000110111010)) color_data = 12'b101001111001;
		if(({row_reg, col_reg}==14'b10000110111011)) color_data = 12'b100101101000;
		if(({row_reg, col_reg}==14'b10000110111100)) color_data = 12'b100001100110;
		if(({row_reg, col_reg}==14'b10000110111101)) color_data = 12'b011101010101;
		if(({row_reg, col_reg}==14'b10000110111110)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==14'b10000110111111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==14'b10000111000000)) color_data = 12'b001100010001;
		if(({row_reg, col_reg}==14'b10000111000001)) color_data = 12'b001100010010;
		if(({row_reg, col_reg}>=14'b10000111000010) && ({row_reg, col_reg}<14'b10000111000100)) color_data = 12'b001100010001;
		if(({row_reg, col_reg}==14'b10000111000100)) color_data = 12'b010100110011;
		if(({row_reg, col_reg}==14'b10000111000101)) color_data = 12'b100101110111;
		if(({row_reg, col_reg}==14'b10000111000110)) color_data = 12'b100101111000;
		if(({row_reg, col_reg}>=14'b10000111000111) && ({row_reg, col_reg}<14'b10000111001001)) color_data = 12'b011101010111;
		if(({row_reg, col_reg}==14'b10000111001001)) color_data = 12'b010100110110;
		if(({row_reg, col_reg}==14'b10000111001010)) color_data = 12'b010100110101;
		if(({row_reg, col_reg}==14'b10000111001011)) color_data = 12'b010101000110;
		if(({row_reg, col_reg}==14'b10000111001100)) color_data = 12'b011101010110;
		if(({row_reg, col_reg}==14'b10000111001101)) color_data = 12'b011001010110;
		if(({row_reg, col_reg}==14'b10000111001110)) color_data = 12'b011101010111;
		if(({row_reg, col_reg}==14'b10000111001111)) color_data = 12'b010100110110;
		if(({row_reg, col_reg}==14'b10000111010000)) color_data = 12'b001000101010;
		if(({row_reg, col_reg}==14'b10000111010001)) color_data = 12'b000100001001;
		if(({row_reg, col_reg}==14'b10000111010010)) color_data = 12'b000000001001;
		if(({row_reg, col_reg}==14'b10000111010011)) color_data = 12'b000000001010;
		if(({row_reg, col_reg}>=14'b10000111010100) && ({row_reg, col_reg}<14'b10000111010110)) color_data = 12'b000000001011;
		if(({row_reg, col_reg}==14'b10000111010110)) color_data = 12'b000000001100;
		if(({row_reg, col_reg}==14'b10000111010111)) color_data = 12'b000000001101;
		if(({row_reg, col_reg}==14'b10000111011000)) color_data = 12'b000000001110;

		if(({row_reg, col_reg}>=14'b10000111011001) && ({row_reg, col_reg}<14'b10001000011100)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==14'b10001000011100)) color_data = 12'b000000001110;
		if(({row_reg, col_reg}==14'b10001000011101)) color_data = 12'b000100001100;
		if(({row_reg, col_reg}==14'b10001000011110)) color_data = 12'b001000001011;
		if(({row_reg, col_reg}==14'b10001000011111)) color_data = 12'b001100001010;
		if(({row_reg, col_reg}>=14'b10001000100000) && ({row_reg, col_reg}<14'b10001000100010)) color_data = 12'b011100010111;
		if(({row_reg, col_reg}==14'b10001000100010)) color_data = 12'b010100000110;
		if(({row_reg, col_reg}==14'b10001000100011)) color_data = 12'b010000000111;
		if(({row_reg, col_reg}==14'b10001000100100)) color_data = 12'b001100001010;
		if(({row_reg, col_reg}==14'b10001000100101)) color_data = 12'b000100001100;
		if(({row_reg, col_reg}>=14'b10001000100110) && ({row_reg, col_reg}<14'b10001000101010)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==14'b10001000101010)) color_data = 12'b000000001100;
		if(({row_reg, col_reg}==14'b10001000101011)) color_data = 12'b000000001010;
		if(({row_reg, col_reg}==14'b10001000101100)) color_data = 12'b000000000111;
		if(({row_reg, col_reg}==14'b10001000101101)) color_data = 12'b000100000110;
		if(({row_reg, col_reg}==14'b10001000101110)) color_data = 12'b000100000101;
		if(({row_reg, col_reg}==14'b10001000101111)) color_data = 12'b001000000100;
		if(({row_reg, col_reg}==14'b10001000110000)) color_data = 12'b001000010011;
		if(({row_reg, col_reg}==14'b10001000110001)) color_data = 12'b001100100011;
		if(({row_reg, col_reg}==14'b10001000110010)) color_data = 12'b011001000101;
		if(({row_reg, col_reg}>=14'b10001000110011) && ({row_reg, col_reg}<14'b10001000110111)) color_data = 12'b011101010110;
		if(({row_reg, col_reg}>=14'b10001000110111) && ({row_reg, col_reg}<14'b10001000111001)) color_data = 12'b100001010111;
		if(({row_reg, col_reg}==14'b10001000111001)) color_data = 12'b100101101000;
		if(({row_reg, col_reg}==14'b10001000111010)) color_data = 12'b100101111000;
		if(({row_reg, col_reg}==14'b10001000111011)) color_data = 12'b101001111000;
		if(({row_reg, col_reg}==14'b10001000111100)) color_data = 12'b101010001000;
		if(({row_reg, col_reg}==14'b10001000111101)) color_data = 12'b100001100110;
		if(({row_reg, col_reg}==14'b10001000111110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==14'b10001000111111)) color_data = 12'b001000000000;
		if(({row_reg, col_reg}==14'b10001001000000)) color_data = 12'b001000000001;
		if(({row_reg, col_reg}==14'b10001001000001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=14'b10001001000010) && ({row_reg, col_reg}<14'b10001001000100)) color_data = 12'b001000000001;
		if(({row_reg, col_reg}==14'b10001001000100)) color_data = 12'b010000100011;
		if(({row_reg, col_reg}>=14'b10001001000101) && ({row_reg, col_reg}<14'b10001001000111)) color_data = 12'b100101111000;
		if(({row_reg, col_reg}==14'b10001001000111)) color_data = 12'b011101010111;
		if(({row_reg, col_reg}==14'b10001001001000)) color_data = 12'b011101011000;
		if(({row_reg, col_reg}==14'b10001001001001)) color_data = 12'b010100110110;
		if(({row_reg, col_reg}==14'b10001001001010)) color_data = 12'b010000100101;
		if(({row_reg, col_reg}==14'b10001001001011)) color_data = 12'b010100110110;
		if(({row_reg, col_reg}==14'b10001001001100)) color_data = 12'b011101010111;
		if(({row_reg, col_reg}>=14'b10001001001101) && ({row_reg, col_reg}<14'b10001001001111)) color_data = 12'b011001000111;
		if(({row_reg, col_reg}==14'b10001001001111)) color_data = 12'b010000100101;
		if(({row_reg, col_reg}==14'b10001001010000)) color_data = 12'b000100011100;
		if(({row_reg, col_reg}==14'b10001001010001)) color_data = 12'b000000001011;
		if(({row_reg, col_reg}==14'b10001001010010)) color_data = 12'b000000001100;
		if(({row_reg, col_reg}==14'b10001001010011)) color_data = 12'b000000001101;
		if(({row_reg, col_reg}>=14'b10001001010100) && ({row_reg, col_reg}<14'b10001001010111)) color_data = 12'b000000001110;

		if(({row_reg, col_reg}>=14'b10001001010111) && ({row_reg, col_reg}<14'b10001010011100)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==14'b10001010011100)) color_data = 12'b000000001110;
		if(({row_reg, col_reg}==14'b10001010011101)) color_data = 12'b000000001101;
		if(({row_reg, col_reg}==14'b10001010011110)) color_data = 12'b001000001011;
		if(({row_reg, col_reg}==14'b10001010011111)) color_data = 12'b001000001010;
		if(({row_reg, col_reg}==14'b10001010100000)) color_data = 12'b001100001010;
		if(({row_reg, col_reg}==14'b10001010100001)) color_data = 12'b010000001010;
		if(({row_reg, col_reg}==14'b10001010100010)) color_data = 12'b001100001001;
		if(({row_reg, col_reg}==14'b10001010100011)) color_data = 12'b001000001010;
		if(({row_reg, col_reg}==14'b10001010100100)) color_data = 12'b000100001100;
		if(({row_reg, col_reg}==14'b10001010100101)) color_data = 12'b000000001110;
		if(({row_reg, col_reg}>=14'b10001010100110) && ({row_reg, col_reg}<14'b10001010101010)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==14'b10001010101010)) color_data = 12'b000000001110;
		if(({row_reg, col_reg}==14'b10001010101011)) color_data = 12'b000000001100;
		if(({row_reg, col_reg}==14'b10001010101100)) color_data = 12'b000000001011;
		if(({row_reg, col_reg}>=14'b10001010101101) && ({row_reg, col_reg}<14'b10001010101111)) color_data = 12'b000000001001;
		if(({row_reg, col_reg}==14'b10001010101111)) color_data = 12'b000100001000;
		if(({row_reg, col_reg}==14'b10001010110000)) color_data = 12'b001000010101;
		if(({row_reg, col_reg}==14'b10001010110001)) color_data = 12'b001000010100;
		if(({row_reg, col_reg}==14'b10001010110010)) color_data = 12'b010000110101;
		if(({row_reg, col_reg}==14'b10001010110011)) color_data = 12'b010100110101;
		if(({row_reg, col_reg}==14'b10001010110100)) color_data = 12'b011001000101;
		if(({row_reg, col_reg}>=14'b10001010110101) && ({row_reg, col_reg}<14'b10001010111001)) color_data = 12'b011101010110;
		if(({row_reg, col_reg}==14'b10001010111001)) color_data = 12'b100101101000;
		if(({row_reg, col_reg}==14'b10001010111010)) color_data = 12'b100001100111;
		if(({row_reg, col_reg}==14'b10001010111011)) color_data = 12'b100101100111;
		if(({row_reg, col_reg}==14'b10001010111100)) color_data = 12'b100101111000;
		if(({row_reg, col_reg}==14'b10001010111101)) color_data = 12'b100101110111;
		if(({row_reg, col_reg}==14'b10001010111110)) color_data = 12'b011101010110;
		if(({row_reg, col_reg}==14'b10001010111111)) color_data = 12'b100001100110;
		if(({row_reg, col_reg}==14'b10001011000000)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==14'b10001011000001)) color_data = 12'b100001100111;
		if(({row_reg, col_reg}==14'b10001011000010)) color_data = 12'b011101010110;
		if(({row_reg, col_reg}==14'b10001011000011)) color_data = 12'b011001000101;
		if(({row_reg, col_reg}==14'b10001011000100)) color_data = 12'b011101010110;
		if(({row_reg, col_reg}==14'b10001011000101)) color_data = 12'b101010001000;
		if(({row_reg, col_reg}==14'b10001011000110)) color_data = 12'b100101111000;
		if(({row_reg, col_reg}==14'b10001011000111)) color_data = 12'b011101010111;
		if(({row_reg, col_reg}==14'b10001011001000)) color_data = 12'b011101011000;
		if(({row_reg, col_reg}==14'b10001011001001)) color_data = 12'b010100110110;
		if(({row_reg, col_reg}==14'b10001011001010)) color_data = 12'b001100010100;
		if(({row_reg, col_reg}==14'b10001011001011)) color_data = 12'b010101000110;
		if(({row_reg, col_reg}>=14'b10001011001100) && ({row_reg, col_reg}<14'b10001011001110)) color_data = 12'b100110001010;
		if(({row_reg, col_reg}==14'b10001011001110)) color_data = 12'b100101111010;
		if(({row_reg, col_reg}==14'b10001011001111)) color_data = 12'b011001000111;
		if(({row_reg, col_reg}==14'b10001011010000)) color_data = 12'b000100011101;
		if(({row_reg, col_reg}==14'b10001011010001)) color_data = 12'b000000001101;
		if(({row_reg, col_reg}==14'b10001011010010)) color_data = 12'b000000001110;

		if(({row_reg, col_reg}>=14'b10001011010011) && ({row_reg, col_reg}<14'b10001100011101)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==14'b10001100011101)) color_data = 12'b000000001110;
		if(({row_reg, col_reg}==14'b10001100011110)) color_data = 12'b000100001101;
		if(({row_reg, col_reg}==14'b10001100011111)) color_data = 12'b000100001100;
		if(({row_reg, col_reg}>=14'b10001100100000) && ({row_reg, col_reg}<14'b10001100100100)) color_data = 12'b000100001101;
		if(({row_reg, col_reg}==14'b10001100100100)) color_data = 12'b000000001110;
		if(({row_reg, col_reg}>=14'b10001100100101) && ({row_reg, col_reg}<14'b10001100101011)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=14'b10001100101011) && ({row_reg, col_reg}<14'b10001100101101)) color_data = 12'b000000001110;
		if(({row_reg, col_reg}>=14'b10001100101101) && ({row_reg, col_reg}<14'b10001100101111)) color_data = 12'b000000001101;
		if(({row_reg, col_reg}==14'b10001100101111)) color_data = 12'b000000001100;
		if(({row_reg, col_reg}==14'b10001100110000)) color_data = 12'b000000000110;
		if(({row_reg, col_reg}==14'b10001100110001)) color_data = 12'b000000000101;
		if(({row_reg, col_reg}==14'b10001100110010)) color_data = 12'b000100000101;
		if(({row_reg, col_reg}==14'b10001100110011)) color_data = 12'b000100000100;
		if(({row_reg, col_reg}==14'b10001100110100)) color_data = 12'b010000100101;
		if(({row_reg, col_reg}==14'b10001100110101)) color_data = 12'b011101010111;
		if(({row_reg, col_reg}>=14'b10001100110110) && ({row_reg, col_reg}<14'b10001100111000)) color_data = 12'b011101010110;
		if(({row_reg, col_reg}==14'b10001100111000)) color_data = 12'b011101010101;
		if(({row_reg, col_reg}==14'b10001100111001)) color_data = 12'b100001010110;
		if(({row_reg, col_reg}==14'b10001100111010)) color_data = 12'b011101010110;
		if(({row_reg, col_reg}==14'b10001100111011)) color_data = 12'b100001100111;
		if(({row_reg, col_reg}==14'b10001100111100)) color_data = 12'b100101110111;
		if(({row_reg, col_reg}==14'b10001100111101)) color_data = 12'b101010001001;
		if(({row_reg, col_reg}==14'b10001100111110)) color_data = 12'b110010101011;
		if(({row_reg, col_reg}==14'b10001100111111)) color_data = 12'b110110111100;
		if(({row_reg, col_reg}==14'b10001101000000)) color_data = 12'b110110111011;
		if(({row_reg, col_reg}==14'b10001101000001)) color_data = 12'b110110111100;
		if(({row_reg, col_reg}==14'b10001101000010)) color_data = 12'b101110011010;
		if(({row_reg, col_reg}==14'b10001101000011)) color_data = 12'b101001111001;
		if(({row_reg, col_reg}>=14'b10001101000100) && ({row_reg, col_reg}<14'b10001101000110)) color_data = 12'b100101111000;
		if(({row_reg, col_reg}>=14'b10001101000110) && ({row_reg, col_reg}<14'b10001101001000)) color_data = 12'b100001100111;
		if(({row_reg, col_reg}==14'b10001101001000)) color_data = 12'b011001000111;
		if(({row_reg, col_reg}==14'b10001101001001)) color_data = 12'b010000100101;
		if(({row_reg, col_reg}==14'b10001101001010)) color_data = 12'b001100010100;
		if(({row_reg, col_reg}==14'b10001101001011)) color_data = 12'b011001010111;
		if(({row_reg, col_reg}==14'b10001101001100)) color_data = 12'b110010111101;
		if(({row_reg, col_reg}==14'b10001101001101)) color_data = 12'b110010101101;
		if(({row_reg, col_reg}==14'b10001101001110)) color_data = 12'b101110101101;
		if(({row_reg, col_reg}==14'b10001101001111)) color_data = 12'b100101111010;
		if(({row_reg, col_reg}==14'b10001101010000)) color_data = 12'b001000101101;
		if(({row_reg, col_reg}==14'b10001101010001)) color_data = 12'b000000001100;
		if(({row_reg, col_reg}==14'b10001101010010)) color_data = 12'b000000001101;

		if(({row_reg, col_reg}>=14'b10001101010011) && ({row_reg, col_reg}<14'b10001110011110)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==14'b10001110011110)) color_data = 12'b000000001110;
		if(({row_reg, col_reg}==14'b10001110011111)) color_data = 12'b000100001110;
		if(({row_reg, col_reg}>=14'b10001110100000) && ({row_reg, col_reg}<14'b10001110101111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==14'b10001110101111)) color_data = 12'b000000001110;
		if(({row_reg, col_reg}==14'b10001110110000)) color_data = 12'b000000001010;
		if(({row_reg, col_reg}==14'b10001110110001)) color_data = 12'b000000001001;
		if(({row_reg, col_reg}==14'b10001110110010)) color_data = 12'b000000001000;
		if(({row_reg, col_reg}==14'b10001110110011)) color_data = 12'b000000000110;
		if(({row_reg, col_reg}==14'b10001110110100)) color_data = 12'b001100100110;
		if(({row_reg, col_reg}==14'b10001110110101)) color_data = 12'b011001010111;
		if(({row_reg, col_reg}>=14'b10001110110110) && ({row_reg, col_reg}<14'b10001110111010)) color_data = 12'b011101010110;
		if(({row_reg, col_reg}==14'b10001110111010)) color_data = 12'b011101000101;
		if(({row_reg, col_reg}>=14'b10001110111011) && ({row_reg, col_reg}<14'b10001110111101)) color_data = 12'b100101111000;
		if(({row_reg, col_reg}==14'b10001110111101)) color_data = 12'b101010001000;
		if(({row_reg, col_reg}==14'b10001110111110)) color_data = 12'b110010011011;
		if(({row_reg, col_reg}==14'b10001110111111)) color_data = 12'b101110011011;
		if(({row_reg, col_reg}==14'b10001111000000)) color_data = 12'b101110011010;
		if(({row_reg, col_reg}==14'b10001111000001)) color_data = 12'b110010101011;
		if(({row_reg, col_reg}==14'b10001111000010)) color_data = 12'b101010001001;
		if(({row_reg, col_reg}==14'b10001111000011)) color_data = 12'b100101111000;
		if(({row_reg, col_reg}==14'b10001111000100)) color_data = 12'b100001100111;
		if(({row_reg, col_reg}==14'b10001111000101)) color_data = 12'b100101111000;
		if(({row_reg, col_reg}==14'b10001111000110)) color_data = 12'b100001100111;
		if(({row_reg, col_reg}==14'b10001111000111)) color_data = 12'b011101010110;
		if(({row_reg, col_reg}==14'b10001111001000)) color_data = 12'b011101010111;
		if(({row_reg, col_reg}==14'b10001111001001)) color_data = 12'b011001000110;
		if(({row_reg, col_reg}==14'b10001111001010)) color_data = 12'b010000110101;
		if(({row_reg, col_reg}==14'b10001111001011)) color_data = 12'b011101100111;
		if(({row_reg, col_reg}==14'b10001111001100)) color_data = 12'b110010111100;
		if(({row_reg, col_reg}>=14'b10001111001101) && ({row_reg, col_reg}<14'b10001111001111)) color_data = 12'b101110101100;
		if(({row_reg, col_reg}==14'b10001111001111)) color_data = 12'b101010011011;
		if(({row_reg, col_reg}==14'b10001111010000)) color_data = 12'b011001011110;
		if(({row_reg, col_reg}==14'b10001111010001)) color_data = 12'b001000101100;
		if(({row_reg, col_reg}==14'b10001111010010)) color_data = 12'b000000001100;
		if(({row_reg, col_reg}==14'b10001111010011)) color_data = 12'b000000001110;

		if(({row_reg, col_reg}>=14'b10001111010100) && ({row_reg, col_reg}<14'b10010000110000)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=14'b10010000110000) && ({row_reg, col_reg}<14'b10010000110010)) color_data = 12'b000000001101;
		if(({row_reg, col_reg}==14'b10010000110010)) color_data = 12'b000000001100;
		if(({row_reg, col_reg}==14'b10010000110011)) color_data = 12'b000100001010;
		if(({row_reg, col_reg}==14'b10010000110100)) color_data = 12'b001100101001;
		if(({row_reg, col_reg}==14'b10010000110101)) color_data = 12'b011101011001;
		if(({row_reg, col_reg}==14'b10010000110110)) color_data = 12'b100101111001;
		if(({row_reg, col_reg}==14'b10010000110111)) color_data = 12'b011101010110;
		if(({row_reg, col_reg}==14'b10010000111000)) color_data = 12'b011101010101;
		if(({row_reg, col_reg}>=14'b10010000111001) && ({row_reg, col_reg}<14'b10010000111011)) color_data = 12'b011101010110;
		if(({row_reg, col_reg}==14'b10010000111011)) color_data = 12'b100001100111;
		if(({row_reg, col_reg}==14'b10010000111100)) color_data = 12'b101001111000;
		if(({row_reg, col_reg}==14'b10010000111101)) color_data = 12'b100101111000;
		if(({row_reg, col_reg}==14'b10010000111110)) color_data = 12'b100101101000;
		if(({row_reg, col_reg}==14'b10010000111111)) color_data = 12'b100101111001;
		if(({row_reg, col_reg}>=14'b10010001000000) && ({row_reg, col_reg}<14'b10010001000011)) color_data = 12'b100101111000;
		if(({row_reg, col_reg}==14'b10010001000011)) color_data = 12'b101010001001;
		if(({row_reg, col_reg}==14'b10010001000100)) color_data = 12'b100001100111;
		if(({row_reg, col_reg}>=14'b10010001000101) && ({row_reg, col_reg}<14'b10010001001000)) color_data = 12'b011101010110;
		if(({row_reg, col_reg}==14'b10010001001000)) color_data = 12'b011001000101;
		if(({row_reg, col_reg}==14'b10010001001001)) color_data = 12'b101010001010;
		if(({row_reg, col_reg}==14'b10010001001010)) color_data = 12'b110010111100;
		if(({row_reg, col_reg}==14'b10010001001011)) color_data = 12'b110010111011;
		if(({row_reg, col_reg}>=14'b10010001001100) && ({row_reg, col_reg}<14'b10010001001110)) color_data = 12'b101110101011;
		if(({row_reg, col_reg}==14'b10010001001110)) color_data = 12'b110010101100;
		if(({row_reg, col_reg}==14'b10010001001111)) color_data = 12'b101110101100;
		if(({row_reg, col_reg}==14'b10010001010000)) color_data = 12'b100110001110;
		if(({row_reg, col_reg}==14'b10010001010001)) color_data = 12'b011001011101;
		if(({row_reg, col_reg}==14'b10010001010010)) color_data = 12'b001100101100;
		if(({row_reg, col_reg}==14'b10010001010011)) color_data = 12'b000000001100;
		if(({row_reg, col_reg}==14'b10010001010100)) color_data = 12'b000000001110;

		if(({row_reg, col_reg}>=14'b10010001010101) && ({row_reg, col_reg}<14'b10010010110010)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==14'b10010010110010)) color_data = 12'b000000001110;
		if(({row_reg, col_reg}==14'b10010010110011)) color_data = 12'b000100001100;
		if(({row_reg, col_reg}==14'b10010010110100)) color_data = 12'b001100101011;
		if(({row_reg, col_reg}==14'b10010010110101)) color_data = 12'b011001011010;
		if(({row_reg, col_reg}==14'b10010010110110)) color_data = 12'b100001111001;
		if(({row_reg, col_reg}==14'b10010010110111)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}>=14'b10010010111000) && ({row_reg, col_reg}<14'b10010010111011)) color_data = 12'b011101010110;
		if(({row_reg, col_reg}==14'b10010010111011)) color_data = 12'b100001100111;
		if(({row_reg, col_reg}==14'b10010010111100)) color_data = 12'b100101111000;
		if(({row_reg, col_reg}==14'b10010010111101)) color_data = 12'b101001111000;
		if(({row_reg, col_reg}==14'b10010010111110)) color_data = 12'b100101111000;
		if(({row_reg, col_reg}==14'b10010010111111)) color_data = 12'b100101111001;
		if(({row_reg, col_reg}==14'b10010011000000)) color_data = 12'b100101111000;
		if(({row_reg, col_reg}>=14'b10010011000001) && ({row_reg, col_reg}<14'b10010011000100)) color_data = 12'b100101111001;
		if(({row_reg, col_reg}==14'b10010011000100)) color_data = 12'b100001100111;
		if(({row_reg, col_reg}>=14'b10010011000101) && ({row_reg, col_reg}<14'b10010011001001)) color_data = 12'b011101010110;
		if(({row_reg, col_reg}==14'b10010011001001)) color_data = 12'b101010001001;
		if(({row_reg, col_reg}>=14'b10010011001010) && ({row_reg, col_reg}<14'b10010011010000)) color_data = 12'b101110101011;
		if(({row_reg, col_reg}==14'b10010011010000)) color_data = 12'b101110101101;
		if(({row_reg, col_reg}==14'b10010011010001)) color_data = 12'b100110001100;
		if(({row_reg, col_reg}==14'b10010011010010)) color_data = 12'b011001011100;
		if(({row_reg, col_reg}==14'b10010011010011)) color_data = 12'b001100101101;
		if(({row_reg, col_reg}==14'b10010011010100)) color_data = 12'b000100001101;

		if(({row_reg, col_reg}>=14'b10010011010101) && ({row_reg, col_reg}<14'b10010100110010)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==14'b10010100110010)) color_data = 12'b000000001110;
		if(({row_reg, col_reg}==14'b10010100110011)) color_data = 12'b000100001101;
		if(({row_reg, col_reg}==14'b10010100110100)) color_data = 12'b001100101011;
		if(({row_reg, col_reg}==14'b10010100110101)) color_data = 12'b011001011010;
		if(({row_reg, col_reg}==14'b10010100110110)) color_data = 12'b100001111001;
		if(({row_reg, col_reg}==14'b10010100110111)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==14'b10010100111000)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}>=14'b10010100111001) && ({row_reg, col_reg}<14'b10010100111011)) color_data = 12'b100101111000;
		if(({row_reg, col_reg}==14'b10010100111011)) color_data = 12'b100101101000;
		if(({row_reg, col_reg}==14'b10010100111100)) color_data = 12'b100001100110;
		if(({row_reg, col_reg}>=14'b10010100111101) && ({row_reg, col_reg}<14'b10010100111111)) color_data = 12'b100001010110;
		if(({row_reg, col_reg}==14'b10010100111111)) color_data = 12'b011101010110;
		if(({row_reg, col_reg}>=14'b10010101000000) && ({row_reg, col_reg}<14'b10010101000010)) color_data = 12'b011101010111;
		if(({row_reg, col_reg}==14'b10010101000010)) color_data = 12'b011001000110;
		if(({row_reg, col_reg}>=14'b10010101000011) && ({row_reg, col_reg}<14'b10010101000101)) color_data = 12'b011000110110;
		if(({row_reg, col_reg}>=14'b10010101000101) && ({row_reg, col_reg}<14'b10010101000111)) color_data = 12'b011101010110;
		if(({row_reg, col_reg}==14'b10010101000111)) color_data = 12'b011001010101;
		if(({row_reg, col_reg}==14'b10010101001000)) color_data = 12'b011001000101;
		if(({row_reg, col_reg}==14'b10010101001001)) color_data = 12'b100001111000;
		if(({row_reg, col_reg}==14'b10010101001010)) color_data = 12'b100110001001;
		if(({row_reg, col_reg}==14'b10010101001011)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==14'b10010101001100)) color_data = 12'b101110101011;
		if(({row_reg, col_reg}==14'b10010101001101)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}>=14'b10010101001110) && ({row_reg, col_reg}<14'b10010101010000)) color_data = 12'b101110101011;
		if(({row_reg, col_reg}==14'b10010101010000)) color_data = 12'b110010111011;
		if(({row_reg, col_reg}==14'b10010101010001)) color_data = 12'b101110101100;
		if(({row_reg, col_reg}==14'b10010101010010)) color_data = 12'b100110001101;
		if(({row_reg, col_reg}==14'b10010101010011)) color_data = 12'b010101011101;
		if(({row_reg, col_reg}==14'b10010101010100)) color_data = 12'b001000101101;
		if(({row_reg, col_reg}==14'b10010101010101)) color_data = 12'b000000001110;

		if(({row_reg, col_reg}>=14'b10010101010110) && ({row_reg, col_reg}<14'b10010110110010)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==14'b10010110110010)) color_data = 12'b000000001110;
		if(({row_reg, col_reg}==14'b10010110110011)) color_data = 12'b001000011100;
		if(({row_reg, col_reg}==14'b10010110110100)) color_data = 12'b010101001011;
		if(({row_reg, col_reg}==14'b10010110110101)) color_data = 12'b011101101010;
		if(({row_reg, col_reg}==14'b10010110110110)) color_data = 12'b100110001001;
		if(({row_reg, col_reg}==14'b10010110110111)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}>=14'b10010110111000) && ({row_reg, col_reg}<14'b10010110111011)) color_data = 12'b100101111000;
		if(({row_reg, col_reg}==14'b10010110111011)) color_data = 12'b100001100111;
		if(({row_reg, col_reg}>=14'b10010110111100) && ({row_reg, col_reg}<14'b10010110111111)) color_data = 12'b011101010110;
		if(({row_reg, col_reg}>=14'b10010110111111) && ({row_reg, col_reg}<14'b10010111000001)) color_data = 12'b011101010111;
		if(({row_reg, col_reg}==14'b10010111000001)) color_data = 12'b100001101000;
		if(({row_reg, col_reg}==14'b10010111000010)) color_data = 12'b010100110110;
		if(({row_reg, col_reg}==14'b10010111000011)) color_data = 12'b010000100101;
		if(({row_reg, col_reg}==14'b10010111000100)) color_data = 12'b010100110110;
		if(({row_reg, col_reg}==14'b10010111000101)) color_data = 12'b011101010111;
		if(({row_reg, col_reg}==14'b10010111000110)) color_data = 12'b011101010110;
		if(({row_reg, col_reg}==14'b10010111000111)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==14'b10010111001000)) color_data = 12'b011001010110;
		if(({row_reg, col_reg}==14'b10010111001001)) color_data = 12'b100001100111;
		if(({row_reg, col_reg}==14'b10010111001010)) color_data = 12'b100001111000;
		if(({row_reg, col_reg}==14'b10010111001011)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==14'b10010111001100)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}>=14'b10010111001101) && ({row_reg, col_reg}<14'b10010111010000)) color_data = 12'b101110101011;
		if(({row_reg, col_reg}==14'b10010111010000)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==14'b10010111010001)) color_data = 12'b101110101011;
		if(({row_reg, col_reg}==14'b10010111010010)) color_data = 12'b101010011101;
		if(({row_reg, col_reg}==14'b10010111010011)) color_data = 12'b100001111110;
		if(({row_reg, col_reg}==14'b10010111010100)) color_data = 12'b010000111110;
		if(({row_reg, col_reg}==14'b10010111010101)) color_data = 12'b000100001101;
		if(({row_reg, col_reg}==14'b10010111010110)) color_data = 12'b000000001110;

		if(({row_reg, col_reg}>=14'b10010111010111) && ({row_reg, col_reg}<14'b10011000110001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==14'b10011000110001)) color_data = 12'b000000001110;
		if(({row_reg, col_reg}==14'b10011000110010)) color_data = 12'b000100011100;
		if(({row_reg, col_reg}==14'b10011000110011)) color_data = 12'b010000111011;
		if(({row_reg, col_reg}==14'b10011000110100)) color_data = 12'b011001101010;
		if(({row_reg, col_reg}==14'b10011000110101)) color_data = 12'b100001111001;
		if(({row_reg, col_reg}>=14'b10011000110110) && ({row_reg, col_reg}<14'b10011000111001)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}>=14'b10011000111001) && ({row_reg, col_reg}<14'b10011000111011)) color_data = 12'b100110001001;
		if(({row_reg, col_reg}==14'b10011000111011)) color_data = 12'b100001100111;
		if(({row_reg, col_reg}>=14'b10011000111100) && ({row_reg, col_reg}<14'b10011000111111)) color_data = 12'b011101010110;
		if(({row_reg, col_reg}==14'b10011000111111)) color_data = 12'b011101010111;
		if(({row_reg, col_reg}==14'b10011001000000)) color_data = 12'b011001010111;
		if(({row_reg, col_reg}==14'b10011001000001)) color_data = 12'b100001101000;
		if(({row_reg, col_reg}==14'b10011001000010)) color_data = 12'b010100110110;
		if(({row_reg, col_reg}==14'b10011001000011)) color_data = 12'b001100010101;
		if(({row_reg, col_reg}==14'b10011001000100)) color_data = 12'b010000100101;
		if(({row_reg, col_reg}==14'b10011001000101)) color_data = 12'b010000100100;
		if(({row_reg, col_reg}==14'b10011001000110)) color_data = 12'b010000100011;
		if(({row_reg, col_reg}==14'b10011001000111)) color_data = 12'b011101100111;
		if(({row_reg, col_reg}==14'b10011001001000)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}>=14'b10011001001001) && ({row_reg, col_reg}<14'b10011001001011)) color_data = 12'b100101111000;
		if(({row_reg, col_reg}==14'b10011001001011)) color_data = 12'b100110001001;
		if(({row_reg, col_reg}==14'b10011001001100)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==14'b10011001001101)) color_data = 12'b101010011010;
		if(({row_reg, col_reg}>=14'b10011001001110) && ({row_reg, col_reg}<14'b10011001010000)) color_data = 12'b101110101011;
		if(({row_reg, col_reg}==14'b10011001010000)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==14'b10011001010001)) color_data = 12'b101110101011;
		if(({row_reg, col_reg}==14'b10011001010010)) color_data = 12'b101110101100;
		if(({row_reg, col_reg}==14'b10011001010011)) color_data = 12'b101010011101;
		if(({row_reg, col_reg}==14'b10011001010100)) color_data = 12'b011001011101;
		if(({row_reg, col_reg}==14'b10011001010101)) color_data = 12'b001000011101;
		if(({row_reg, col_reg}==14'b10011001010110)) color_data = 12'b000000001101;

		if(({row_reg, col_reg}>=14'b10011001010111) && ({row_reg, col_reg}<14'b10011010110000)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==14'b10011010110000)) color_data = 12'b000000001110;
		if(({row_reg, col_reg}==14'b10011010110001)) color_data = 12'b000000001101;
		if(({row_reg, col_reg}==14'b10011010110010)) color_data = 12'b001000101011;
		if(({row_reg, col_reg}==14'b10011010110011)) color_data = 12'b010101011010;
		if(({row_reg, col_reg}==14'b10011010110100)) color_data = 12'b011101111001;
		if(({row_reg, col_reg}==14'b10011010110101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=14'b10011010110110) && ({row_reg, col_reg}<14'b10011010111001)) color_data = 12'b100101111000;
		if(({row_reg, col_reg}==14'b10011010111001)) color_data = 12'b100110001001;
		if(({row_reg, col_reg}==14'b10011010111010)) color_data = 12'b101010001001;
		if(({row_reg, col_reg}==14'b10011010111011)) color_data = 12'b100001111000;
		if(({row_reg, col_reg}==14'b10011010111100)) color_data = 12'b011101010111;
		if(({row_reg, col_reg}==14'b10011010111101)) color_data = 12'b011101100111;
		if(({row_reg, col_reg}>=14'b10011010111110) && ({row_reg, col_reg}<14'b10011011000001)) color_data = 12'b011101010111;
		if(({row_reg, col_reg}==14'b10011011000001)) color_data = 12'b011101011000;
		if(({row_reg, col_reg}==14'b10011011000010)) color_data = 12'b010100110110;
		if(({row_reg, col_reg}>=14'b10011011000011) && ({row_reg, col_reg}<14'b10011011000101)) color_data = 12'b001100010100;
		if(({row_reg, col_reg}>=14'b10011011000101) && ({row_reg, col_reg}<14'b10011011000111)) color_data = 12'b001100010010;
		if(({row_reg, col_reg}==14'b10011011000111)) color_data = 12'b100101111000;
		if(({row_reg, col_reg}>=14'b10011011001000) && ({row_reg, col_reg}<14'b10011011001100)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==14'b10011011001100)) color_data = 12'b100001111000;
		if(({row_reg, col_reg}==14'b10011011001101)) color_data = 12'b100110001001;
		if(({row_reg, col_reg}==14'b10011011001110)) color_data = 12'b101110101011;
		if(({row_reg, col_reg}==14'b10011011001111)) color_data = 12'b110010101011;
		if(({row_reg, col_reg}==14'b10011011010000)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}>=14'b10011011010001) && ({row_reg, col_reg}<14'b10011011010011)) color_data = 12'b101110101011;
		if(({row_reg, col_reg}==14'b10011011010011)) color_data = 12'b101110101100;
		if(({row_reg, col_reg}==14'b10011011010100)) color_data = 12'b100001111100;
		if(({row_reg, col_reg}==14'b10011011010101)) color_data = 12'b010000111100;
		if(({row_reg, col_reg}==14'b10011011010110)) color_data = 12'b000100001100;
		if(({row_reg, col_reg}==14'b10011011010111)) color_data = 12'b000000001101;

		if(({row_reg, col_reg}>=14'b10011011011000) && ({row_reg, col_reg}<14'b10011100110000)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==14'b10011100110000)) color_data = 12'b000000001110;
		if(({row_reg, col_reg}==14'b10011100110001)) color_data = 12'b000100001100;
		if(({row_reg, col_reg}==14'b10011100110010)) color_data = 12'b010001001100;
		if(({row_reg, col_reg}==14'b10011100110011)) color_data = 12'b100001111011;
		if(({row_reg, col_reg}==14'b10011100110100)) color_data = 12'b100110001010;
		if(({row_reg, col_reg}==14'b10011100110101)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}>=14'b10011100110110) && ({row_reg, col_reg}<14'b10011100111000)) color_data = 12'b101010001001;
		if(({row_reg, col_reg}==14'b10011100111000)) color_data = 12'b101010001010;
		if(({row_reg, col_reg}>=14'b10011100111001) && ({row_reg, col_reg}<14'b10011100111011)) color_data = 12'b100001111000;
		if(({row_reg, col_reg}==14'b10011100111011)) color_data = 12'b011101100111;
		if(({row_reg, col_reg}>=14'b10011100111100) && ({row_reg, col_reg}<14'b10011100111111)) color_data = 12'b011001000110;
		if(({row_reg, col_reg}==14'b10011100111111)) color_data = 12'b011001000111;
		if(({row_reg, col_reg}==14'b10011101000000)) color_data = 12'b011001010111;
		if(({row_reg, col_reg}==14'b10011101000001)) color_data = 12'b011001000111;
		if(({row_reg, col_reg}==14'b10011101000010)) color_data = 12'b010000100101;
		if(({row_reg, col_reg}==14'b10011101000011)) color_data = 12'b001100010100;
		if(({row_reg, col_reg}==14'b10011101000100)) color_data = 12'b001100010011;
		if(({row_reg, col_reg}==14'b10011101000101)) color_data = 12'b001100010010;
		if(({row_reg, col_reg}==14'b10011101000110)) color_data = 12'b001100010001;
		if(({row_reg, col_reg}==14'b10011101000111)) color_data = 12'b100101111000;
		if(({row_reg, col_reg}>=14'b10011101001000) && ({row_reg, col_reg}<14'b10011101001100)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==14'b10011101001100)) color_data = 12'b100101111000;
		if(({row_reg, col_reg}==14'b10011101001101)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==14'b10011101001110)) color_data = 12'b101110011010;
		if(({row_reg, col_reg}==14'b10011101001111)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==14'b10011101010000)) color_data = 12'b101110101011;
		if(({row_reg, col_reg}==14'b10011101010001)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==14'b10011101010010)) color_data = 12'b101110111010;
		if(({row_reg, col_reg}==14'b10011101010011)) color_data = 12'b101110101011;
		if(({row_reg, col_reg}==14'b10011101010100)) color_data = 12'b101010011100;
		if(({row_reg, col_reg}==14'b10011101010101)) color_data = 12'b011001101100;
		if(({row_reg, col_reg}==14'b10011101010110)) color_data = 12'b001100101100;
		if(({row_reg, col_reg}==14'b10011101010111)) color_data = 12'b000000001101;
		if(({row_reg, col_reg}==14'b10011101011000)) color_data = 12'b000000001110;

		if(({row_reg, col_reg}>=14'b10011101011001) && ({row_reg, col_reg}<14'b10011110110001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==14'b10011110110001)) color_data = 12'b001000011101;
		if(({row_reg, col_reg}==14'b10011110110010)) color_data = 12'b011001101101;
		if(({row_reg, col_reg}==14'b10011110110011)) color_data = 12'b101010101100;
		if(({row_reg, col_reg}==14'b10011110110100)) color_data = 12'b101110101011;
		if(({row_reg, col_reg}==14'b10011110110101)) color_data = 12'b110010111011;
		if(({row_reg, col_reg}==14'b10011110110110)) color_data = 12'b110010101011;
		if(({row_reg, col_reg}==14'b10011110110111)) color_data = 12'b110010101100;
		if(({row_reg, col_reg}==14'b10011110111000)) color_data = 12'b110010111101;
		if(({row_reg, col_reg}==14'b10011110111001)) color_data = 12'b011101010111;
		if(({row_reg, col_reg}>=14'b10011110111010) && ({row_reg, col_reg}<14'b10011110111100)) color_data = 12'b010100110101;
		if(({row_reg, col_reg}==14'b10011110111100)) color_data = 12'b010000100100;
		if(({row_reg, col_reg}>=14'b10011110111101) && ({row_reg, col_reg}<14'b10011111000000)) color_data = 12'b010000100101;
		if(({row_reg, col_reg}>=14'b10011111000000) && ({row_reg, col_reg}<14'b10011111000011)) color_data = 12'b010000100100;
		if(({row_reg, col_reg}==14'b10011111000011)) color_data = 12'b001000010011;
		if(({row_reg, col_reg}==14'b10011111000100)) color_data = 12'b001100010011;
		if(({row_reg, col_reg}==14'b10011111000101)) color_data = 12'b001100010010;
		if(({row_reg, col_reg}==14'b10011111000110)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==14'b10011111000111)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}>=14'b10011111001000) && ({row_reg, col_reg}<14'b10011111001010)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==14'b10011111001010)) color_data = 12'b100101111000;
		if(({row_reg, col_reg}>=14'b10011111001011) && ({row_reg, col_reg}<14'b10011111001101)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}>=14'b10011111001101) && ({row_reg, col_reg}<14'b10011111010000)) color_data = 12'b100101111000;
		if(({row_reg, col_reg}>=14'b10011111010000) && ({row_reg, col_reg}<14'b10011111010010)) color_data = 12'b101110101011;
		if(({row_reg, col_reg}>=14'b10011111010010) && ({row_reg, col_reg}<14'b10011111010100)) color_data = 12'b101110111010;
		if(({row_reg, col_reg}==14'b10011111010100)) color_data = 12'b101110101100;
		if(({row_reg, col_reg}==14'b10011111010101)) color_data = 12'b100110001101;
		if(({row_reg, col_reg}==14'b10011111010110)) color_data = 12'b010101011101;
		if(({row_reg, col_reg}==14'b10011111010111)) color_data = 12'b001000101101;
		if(({row_reg, col_reg}==14'b10011111011000)) color_data = 12'b000000001110;

		if(({row_reg, col_reg}>=14'b10011111011001) && ({row_reg, col_reg}<14'b10100000101111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==14'b10100000101111)) color_data = 12'b000000001110;
		if(({row_reg, col_reg}==14'b10100000110000)) color_data = 12'b000100001100;
		if(({row_reg, col_reg}==14'b10100000110001)) color_data = 12'b010101001101;
		if(({row_reg, col_reg}==14'b10100000110010)) color_data = 12'b100010001100;
		if(({row_reg, col_reg}==14'b10100000110011)) color_data = 12'b101110101100;
		if(({row_reg, col_reg}==14'b10100000110100)) color_data = 12'b110010101011;
		if(({row_reg, col_reg}==14'b10100000110101)) color_data = 12'b101110011011;
		if(({row_reg, col_reg}==14'b10100000110110)) color_data = 12'b110010101100;
		if(({row_reg, col_reg}==14'b10100000110111)) color_data = 12'b101110011100;
		if(({row_reg, col_reg}==14'b10100000111000)) color_data = 12'b101110101100;
		if(({row_reg, col_reg}==14'b10100000111001)) color_data = 12'b011101011000;
		if(({row_reg, col_reg}>=14'b10100000111010) && ({row_reg, col_reg}<14'b10100000111100)) color_data = 12'b010100110111;
		if(({row_reg, col_reg}==14'b10100000111100)) color_data = 12'b010000100110;
		if(({row_reg, col_reg}>=14'b10100000111101) && ({row_reg, col_reg}<14'b10100001000000)) color_data = 12'b010000100101;
		if(({row_reg, col_reg}==14'b10100001000000)) color_data = 12'b010000110100;
		if(({row_reg, col_reg}==14'b10100001000001)) color_data = 12'b010100110100;
		if(({row_reg, col_reg}==14'b10100001000010)) color_data = 12'b001100100011;
		if(({row_reg, col_reg}>=14'b10100001000011) && ({row_reg, col_reg}<14'b10100001000101)) color_data = 12'b001100010010;
		if(({row_reg, col_reg}==14'b10100001000101)) color_data = 12'b001100010001;
		if(({row_reg, col_reg}==14'b10100001000110)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}==14'b10100001000111)) color_data = 12'b100001100111;
		if(({row_reg, col_reg}>=14'b10100001001000) && ({row_reg, col_reg}<14'b10100001001010)) color_data = 12'b100101111000;
		if(({row_reg, col_reg}==14'b10100001001010)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==14'b10100001001011)) color_data = 12'b100101110111;
		if(({row_reg, col_reg}>=14'b10100001001100) && ({row_reg, col_reg}<14'b10100001010000)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==14'b10100001010000)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==14'b10100001010001)) color_data = 12'b101110101011;
		if(({row_reg, col_reg}>=14'b10100001010010) && ({row_reg, col_reg}<14'b10100001010100)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==14'b10100001010100)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==14'b10100001010101)) color_data = 12'b101110101011;
		if(({row_reg, col_reg}==14'b10100001010110)) color_data = 12'b100110001100;
		if(({row_reg, col_reg}==14'b10100001010111)) color_data = 12'b010101001011;
		if(({row_reg, col_reg}==14'b10100001011000)) color_data = 12'b001000011100;
		if(({row_reg, col_reg}==14'b10100001011001)) color_data = 12'b000000001101;

		if(({row_reg, col_reg}>=14'b10100001011010) && ({row_reg, col_reg}<14'b10100010110000)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==14'b10100010110000)) color_data = 12'b001000011101;
		if(({row_reg, col_reg}==14'b10100010110001)) color_data = 12'b011001101110;
		if(({row_reg, col_reg}==14'b10100010110010)) color_data = 12'b101010011110;
		if(({row_reg, col_reg}==14'b10100010110011)) color_data = 12'b110010111100;
		if(({row_reg, col_reg}==14'b10100010110100)) color_data = 12'b100110001001;
		if(({row_reg, col_reg}>=14'b10100010110101) && ({row_reg, col_reg}<14'b10100010110111)) color_data = 12'b011001000110;
		if(({row_reg, col_reg}>=14'b10100010110111) && ({row_reg, col_reg}<14'b10100010111001)) color_data = 12'b011001000111;
		if(({row_reg, col_reg}==14'b10100010111001)) color_data = 12'b010101000111;
		if(({row_reg, col_reg}==14'b10100010111010)) color_data = 12'b011001000111;
		if(({row_reg, col_reg}==14'b10100010111011)) color_data = 12'b010100110111;
		if(({row_reg, col_reg}==14'b10100010111100)) color_data = 12'b010000100101;
		if(({row_reg, col_reg}>=14'b10100010111101) && ({row_reg, col_reg}<14'b10100011000000)) color_data = 12'b010000110101;
		if(({row_reg, col_reg}==14'b10100011000000)) color_data = 12'b100001101000;
		if(({row_reg, col_reg}==14'b10100011000001)) color_data = 12'b100110001001;
		if(({row_reg, col_reg}==14'b10100011000010)) color_data = 12'b010101000101;
		if(({row_reg, col_reg}==14'b10100011000011)) color_data = 12'b001000000001;
		if(({row_reg, col_reg}>=14'b10100011000100) && ({row_reg, col_reg}<14'b10100011000110)) color_data = 12'b001100010010;
		if(({row_reg, col_reg}==14'b10100011000110)) color_data = 12'b001100010001;
		if(({row_reg, col_reg}==14'b10100011000111)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}==14'b10100011001000)) color_data = 12'b001100010001;
		if(({row_reg, col_reg}==14'b10100011001001)) color_data = 12'b011101010110;
		if(({row_reg, col_reg}>=14'b10100011001010) && ({row_reg, col_reg}<14'b10100011001100)) color_data = 12'b101010001000;
		if(({row_reg, col_reg}>=14'b10100011001100) && ({row_reg, col_reg}<14'b10100011010010)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==14'b10100011010010)) color_data = 12'b101010011010;
		if(({row_reg, col_reg}>=14'b10100011010011) && ({row_reg, col_reg}<14'b10100011010101)) color_data = 12'b110010111011;
		if(({row_reg, col_reg}==14'b10100011010101)) color_data = 12'b101110101011;
		if(({row_reg, col_reg}==14'b10100011010110)) color_data = 12'b101110101100;
		if(({row_reg, col_reg}==14'b10100011010111)) color_data = 12'b100001111101;
		if(({row_reg, col_reg}==14'b10100011011000)) color_data = 12'b010001001101;
		if(({row_reg, col_reg}==14'b10100011011001)) color_data = 12'b000100011101;
		if(({row_reg, col_reg}==14'b10100011011010)) color_data = 12'b000000001110;

		if(({row_reg, col_reg}>=14'b10100011011011) && ({row_reg, col_reg}<14'b10100100101111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==14'b10100100101111)) color_data = 12'b000000001110;
		if(({row_reg, col_reg}==14'b10100100110000)) color_data = 12'b010001001101;
		if(({row_reg, col_reg}==14'b10100100110001)) color_data = 12'b100001111110;
		if(({row_reg, col_reg}==14'b10100100110010)) color_data = 12'b101110101110;
		if(({row_reg, col_reg}==14'b10100100110011)) color_data = 12'b110010111101;
		if(({row_reg, col_reg}==14'b10100100110100)) color_data = 12'b100101111001;
		if(({row_reg, col_reg}>=14'b10100100110101) && ({row_reg, col_reg}<14'b10100100110111)) color_data = 12'b010100110110;
		if(({row_reg, col_reg}==14'b10100100110111)) color_data = 12'b011001000111;
		if(({row_reg, col_reg}==14'b10100100111000)) color_data = 12'b010100110110;
		if(({row_reg, col_reg}==14'b10100100111001)) color_data = 12'b011001000111;
		if(({row_reg, col_reg}==14'b10100100111010)) color_data = 12'b011001001000;
		if(({row_reg, col_reg}==14'b10100100111011)) color_data = 12'b010000110110;
		if(({row_reg, col_reg}>=14'b10100100111100) && ({row_reg, col_reg}<14'b10100100111110)) color_data = 12'b001100100100;
		if(({row_reg, col_reg}==14'b10100100111110)) color_data = 12'b001100010011;
		if(({row_reg, col_reg}==14'b10100100111111)) color_data = 12'b001100100100;
		if(({row_reg, col_reg}==14'b10100101000000)) color_data = 12'b100001111000;
		if(({row_reg, col_reg}==14'b10100101000001)) color_data = 12'b101010001001;
		if(({row_reg, col_reg}==14'b10100101000010)) color_data = 12'b011001000101;
		if(({row_reg, col_reg}==14'b10100101000011)) color_data = 12'b001000000001;
		if(({row_reg, col_reg}==14'b10100101000100)) color_data = 12'b001100010001;
		if(({row_reg, col_reg}==14'b10100101000101)) color_data = 12'b001100010010;
		if(({row_reg, col_reg}>=14'b10100101000110) && ({row_reg, col_reg}<14'b10100101001000)) color_data = 12'b001100010001;
		if(({row_reg, col_reg}==14'b10100101001000)) color_data = 12'b001000000000;
		if(({row_reg, col_reg}==14'b10100101001001)) color_data = 12'b011101010101;
		if(({row_reg, col_reg}>=14'b10100101001010) && ({row_reg, col_reg}<14'b10100101001100)) color_data = 12'b101010001000;
		if(({row_reg, col_reg}>=14'b10100101001100) && ({row_reg, col_reg}<14'b10100101001110)) color_data = 12'b100101111000;
		if(({row_reg, col_reg}==14'b10100101001110)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==14'b10100101001111)) color_data = 12'b100101111000;
		if(({row_reg, col_reg}==14'b10100101010000)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==14'b10100101010001)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==14'b10100101010010)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==14'b10100101010011)) color_data = 12'b101110101011;
		if(({row_reg, col_reg}==14'b10100101010100)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==14'b10100101010101)) color_data = 12'b101110101011;
		if(({row_reg, col_reg}==14'b10100101010110)) color_data = 12'b101110101100;
		if(({row_reg, col_reg}==14'b10100101010111)) color_data = 12'b101010011101;
		if(({row_reg, col_reg}==14'b10100101011000)) color_data = 12'b011101101110;
		if(({row_reg, col_reg}==14'b10100101011001)) color_data = 12'b001100111101;
		if(({row_reg, col_reg}==14'b10100101011010)) color_data = 12'b000000001101;
		if(({row_reg, col_reg}==14'b10100101011011)) color_data = 12'b000000001110;

		if(({row_reg, col_reg}>=14'b10100101011100) && ({row_reg, col_reg}<14'b10100110101110)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=14'b10100110101110) && ({row_reg, col_reg}<14'b10100110110000)) color_data = 12'b000000001110;
		if(({row_reg, col_reg}==14'b10100110110000)) color_data = 12'b001100111010;
		if(({row_reg, col_reg}==14'b10100110110001)) color_data = 12'b011001011011;
		if(({row_reg, col_reg}==14'b10100110110010)) color_data = 12'b011101101010;
		if(({row_reg, col_reg}==14'b10100110110011)) color_data = 12'b100001101001;
		if(({row_reg, col_reg}==14'b10100110110100)) color_data = 12'b011101011000;
		if(({row_reg, col_reg}==14'b10100110110101)) color_data = 12'b011001000111;
		if(({row_reg, col_reg}==14'b10100110110110)) color_data = 12'b011001001000;
		if(({row_reg, col_reg}==14'b10100110110111)) color_data = 12'b010101000111;
		if(({row_reg, col_reg}==14'b10100110111000)) color_data = 12'b011001001000;
		if(({row_reg, col_reg}==14'b10100110111001)) color_data = 12'b010000110110;
		if(({row_reg, col_reg}==14'b10100110111010)) color_data = 12'b010000100110;
		if(({row_reg, col_reg}==14'b10100110111011)) color_data = 12'b011101011000;
		if(({row_reg, col_reg}==14'b10100110111100)) color_data = 12'b101010001010;
		if(({row_reg, col_reg}==14'b10100110111101)) color_data = 12'b100110001001;
		if(({row_reg, col_reg}==14'b10100110111110)) color_data = 12'b011101100111;
		if(({row_reg, col_reg}>=14'b10100110111111) && ({row_reg, col_reg}<14'b10100111000001)) color_data = 12'b100001111000;
		if(({row_reg, col_reg}==14'b10100111000001)) color_data = 12'b100110001001;
		if(({row_reg, col_reg}==14'b10100111000010)) color_data = 12'b010101000101;
		if(({row_reg, col_reg}==14'b10100111000011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==14'b10100111000100)) color_data = 12'b001100010010;
		if(({row_reg, col_reg}>=14'b10100111000101) && ({row_reg, col_reg}<14'b10100111001001)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}==14'b10100111001001)) color_data = 12'b010100110011;
		if(({row_reg, col_reg}>=14'b10100111001010) && ({row_reg, col_reg}<14'b10100111001100)) color_data = 12'b010100110100;
		if(({row_reg, col_reg}==14'b10100111001100)) color_data = 12'b010100110011;
		if(({row_reg, col_reg}==14'b10100111001101)) color_data = 12'b011001000100;
		if(({row_reg, col_reg}==14'b10100111001110)) color_data = 12'b100101110111;
		if(({row_reg, col_reg}==14'b10100111001111)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==14'b10100111010000)) color_data = 12'b101010001001;
		if(({row_reg, col_reg}==14'b10100111010001)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==14'b10100111010010)) color_data = 12'b101010001001;
		if(({row_reg, col_reg}==14'b10100111010011)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==14'b10100111010100)) color_data = 12'b101010011000;
		if(({row_reg, col_reg}==14'b10100111010101)) color_data = 12'b101110111010;
		if(({row_reg, col_reg}==14'b10100111010110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==14'b10100111010111)) color_data = 12'b101110101100;
		if(({row_reg, col_reg}==14'b10100111011000)) color_data = 12'b100110001101;
		if(({row_reg, col_reg}==14'b10100111011001)) color_data = 12'b010101011101;
		if(({row_reg, col_reg}==14'b10100111011010)) color_data = 12'b000100011100;
		if(({row_reg, col_reg}==14'b10100111011011)) color_data = 12'b000000001101;

		if(({row_reg, col_reg}>=14'b10100111011100) && ({row_reg, col_reg}<14'b10101000101110)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==14'b10101000101110)) color_data = 12'b000000001101;
		if(({row_reg, col_reg}==14'b10101000101111)) color_data = 12'b000100011101;
		if(({row_reg, col_reg}==14'b10101000110000)) color_data = 12'b001100101000;
		if(({row_reg, col_reg}==14'b10101000110001)) color_data = 12'b010000111000;
		if(({row_reg, col_reg}==14'b10101000110010)) color_data = 12'b010000110110;
		if(({row_reg, col_reg}>=14'b10101000110011) && ({row_reg, col_reg}<14'b10101000110101)) color_data = 12'b010100110110;
		if(({row_reg, col_reg}==14'b10101000110101)) color_data = 12'b010100110111;
		if(({row_reg, col_reg}==14'b10101000110110)) color_data = 12'b011001001000;
		if(({row_reg, col_reg}==14'b10101000110111)) color_data = 12'b010100110111;
		if(({row_reg, col_reg}==14'b10101000111000)) color_data = 12'b011001000111;
		if(({row_reg, col_reg}==14'b10101000111001)) color_data = 12'b010000100101;
		if(({row_reg, col_reg}==14'b10101000111010)) color_data = 12'b001100010100;
		if(({row_reg, col_reg}==14'b10101000111011)) color_data = 12'b011101101000;
		if(({row_reg, col_reg}==14'b10101000111100)) color_data = 12'b110110111101;
		if(({row_reg, col_reg}==14'b10101000111101)) color_data = 12'b110010101011;
		if(({row_reg, col_reg}==14'b10101000111110)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==14'b10101000111111)) color_data = 12'b100110001001;
		if(({row_reg, col_reg}==14'b10101001000000)) color_data = 12'b101010001001;
		if(({row_reg, col_reg}==14'b10101001000001)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==14'b10101001000010)) color_data = 12'b011001000101;
		if(({row_reg, col_reg}==14'b10101001000011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==14'b10101001000100)) color_data = 12'b001100010001;
		if(({row_reg, col_reg}>=14'b10101001000101) && ({row_reg, col_reg}<14'b10101001000111)) color_data = 12'b010100110011;
		if(({row_reg, col_reg}>=14'b10101001000111) && ({row_reg, col_reg}<14'b10101001001001)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}==14'b10101001001001)) color_data = 12'b001100010001;
		if(({row_reg, col_reg}>=14'b10101001001010) && ({row_reg, col_reg}<14'b10101001001101)) color_data = 12'b001000000000;
		if(({row_reg, col_reg}==14'b10101001001101)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}==14'b10101001001110)) color_data = 12'b100101110111;
		if(({row_reg, col_reg}==14'b10101001001111)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}>=14'b10101001010000) && ({row_reg, col_reg}<14'b10101001010101)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==14'b10101001010101)) color_data = 12'b110010111010;
		if(({row_reg, col_reg}==14'b10101001010110)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==14'b10101001010111)) color_data = 12'b101110111100;
		if(({row_reg, col_reg}==14'b10101001011000)) color_data = 12'b101010011101;
		if(({row_reg, col_reg}==14'b10101001011001)) color_data = 12'b011101111101;
		if(({row_reg, col_reg}==14'b10101001011010)) color_data = 12'b001100111101;
		if(({row_reg, col_reg}==14'b10101001011011)) color_data = 12'b000000001100;
		if(({row_reg, col_reg}==14'b10101001011100)) color_data = 12'b000000001110;

		if(({row_reg, col_reg}>=14'b10101001011101) && ({row_reg, col_reg}<14'b10101010101101)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==14'b10101010101101)) color_data = 12'b000000001101;
		if(({row_reg, col_reg}==14'b10101010101110)) color_data = 12'b000000001100;
		if(({row_reg, col_reg}==14'b10101010101111)) color_data = 12'b001000011011;
		if(({row_reg, col_reg}==14'b10101010110000)) color_data = 12'b010000111000;
		if(({row_reg, col_reg}==14'b10101010110001)) color_data = 12'b010101001000;
		if(({row_reg, col_reg}==14'b10101010110010)) color_data = 12'b010101000111;
		if(({row_reg, col_reg}==14'b10101010110011)) color_data = 12'b011001000111;
		if(({row_reg, col_reg}==14'b10101010110100)) color_data = 12'b010101000111;
		if(({row_reg, col_reg}>=14'b10101010110101) && ({row_reg, col_reg}<14'b10101010111000)) color_data = 12'b010100110111;
		if(({row_reg, col_reg}==14'b10101010111000)) color_data = 12'b010000110110;
		if(({row_reg, col_reg}==14'b10101010111001)) color_data = 12'b011001011000;
		if(({row_reg, col_reg}==14'b10101010111010)) color_data = 12'b011101011000;
		if(({row_reg, col_reg}==14'b10101010111011)) color_data = 12'b100101111001;
		if(({row_reg, col_reg}==14'b10101010111100)) color_data = 12'b110010111011;
		if(({row_reg, col_reg}==14'b10101010111101)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==14'b10101010111110)) color_data = 12'b100001111000;
		if(({row_reg, col_reg}==14'b10101010111111)) color_data = 12'b100110001001;
		if(({row_reg, col_reg}>=14'b10101011000000) && ({row_reg, col_reg}<14'b10101011000010)) color_data = 12'b011101010110;
		if(({row_reg, col_reg}==14'b10101011000010)) color_data = 12'b010000110011;
		if(({row_reg, col_reg}==14'b10101011000011)) color_data = 12'b001000000001;
		if(({row_reg, col_reg}==14'b10101011000100)) color_data = 12'b001100010001;
		if(({row_reg, col_reg}==14'b10101011000101)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==14'b10101011000110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==14'b10101011000111)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}==14'b10101011001000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==14'b10101011001001)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}==14'b10101011001010)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==14'b10101011001011)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}==14'b10101011001100)) color_data = 12'b001100010001;
		if(({row_reg, col_reg}==14'b10101011001101)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}==14'b10101011001110)) color_data = 12'b011001010101;
		if(({row_reg, col_reg}==14'b10101011001111)) color_data = 12'b011101010101;
		if(({row_reg, col_reg}==14'b10101011010000)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==14'b10101011010001)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==14'b10101011010010)) color_data = 12'b100101111000;
		if(({row_reg, col_reg}>=14'b10101011010011) && ({row_reg, col_reg}<14'b10101011010101)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==14'b10101011010101)) color_data = 12'b101110011001;
		if(({row_reg, col_reg}==14'b10101011010110)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==14'b10101011010111)) color_data = 12'b101110101011;
		if(({row_reg, col_reg}==14'b10101011011000)) color_data = 12'b101110101100;
		if(({row_reg, col_reg}==14'b10101011011001)) color_data = 12'b101010011101;
		if(({row_reg, col_reg}==14'b10101011011010)) color_data = 12'b011001101101;
		if(({row_reg, col_reg}==14'b10101011011011)) color_data = 12'b001000101101;
		if(({row_reg, col_reg}==14'b10101011011100)) color_data = 12'b000000001101;

		if(({row_reg, col_reg}>=14'b10101011011101) && ({row_reg, col_reg}<14'b10101100101011)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=14'b10101100101011) && ({row_reg, col_reg}<14'b10101100101101)) color_data = 12'b000000001110;
		if(({row_reg, col_reg}==14'b10101100101101)) color_data = 12'b000000001100;
		if(({row_reg, col_reg}==14'b10101100101110)) color_data = 12'b000100001010;
		if(({row_reg, col_reg}==14'b10101100101111)) color_data = 12'b001100101001;
		if(({row_reg, col_reg}==14'b10101100110000)) color_data = 12'b010000111000;
		if(({row_reg, col_reg}==14'b10101100110001)) color_data = 12'b010101001000;
		if(({row_reg, col_reg}==14'b10101100110010)) color_data = 12'b010101000111;
		if(({row_reg, col_reg}==14'b10101100110011)) color_data = 12'b011001000111;
		if(({row_reg, col_reg}==14'b10101100110100)) color_data = 12'b010100110110;
		if(({row_reg, col_reg}>=14'b10101100110101) && ({row_reg, col_reg}<14'b10101100111000)) color_data = 12'b001100100101;
		if(({row_reg, col_reg}==14'b10101100111000)) color_data = 12'b001100100100;
		if(({row_reg, col_reg}==14'b10101100111001)) color_data = 12'b100110001010;
		if(({row_reg, col_reg}==14'b10101100111010)) color_data = 12'b110010101100;
		if(({row_reg, col_reg}==14'b10101100111011)) color_data = 12'b110010101011;
		if(({row_reg, col_reg}==14'b10101100111100)) color_data = 12'b110010111011;
		if(({row_reg, col_reg}==14'b10101100111101)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}>=14'b10101100111110) && ({row_reg, col_reg}<14'b10101101000000)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==14'b10101101000000)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}>=14'b10101101000001) && ({row_reg, col_reg}<14'b10101101000100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==14'b10101101000100)) color_data = 12'b001100010001;
		if(({row_reg, col_reg}>=14'b10101101000101) && ({row_reg, col_reg}<14'b10101101000111)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}==14'b10101101000111)) color_data = 12'b010100110011;
		if(({row_reg, col_reg}>=14'b10101101001000) && ({row_reg, col_reg}<14'b10101101001010)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}==14'b10101101001010)) color_data = 12'b010000100011;
		if(({row_reg, col_reg}==14'b10101101001011)) color_data = 12'b010000110011;
		if(({row_reg, col_reg}>=14'b10101101001100) && ({row_reg, col_reg}<14'b10101101001110)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}==14'b10101101001110)) color_data = 12'b001100010001;
		if(({row_reg, col_reg}==14'b10101101001111)) color_data = 12'b001000000000;
		if(({row_reg, col_reg}==14'b10101101010000)) color_data = 12'b100001100110;
		if(({row_reg, col_reg}==14'b10101101010001)) color_data = 12'b101010001000;
		if(({row_reg, col_reg}==14'b10101101010010)) color_data = 12'b100101111000;
		if(({row_reg, col_reg}>=14'b10101101010011) && ({row_reg, col_reg}<14'b10101101010110)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==14'b10101101010110)) color_data = 12'b100110000111;
		if(({row_reg, col_reg}==14'b10101101010111)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==14'b10101101011000)) color_data = 12'b101110101011;
		if(({row_reg, col_reg}==14'b10101101011001)) color_data = 12'b101110101101;
		if(({row_reg, col_reg}==14'b10101101011010)) color_data = 12'b100110001110;
		if(({row_reg, col_reg}==14'b10101101011011)) color_data = 12'b010101001101;
		if(({row_reg, col_reg}==14'b10101101011100)) color_data = 12'b000100011101;
		if(({row_reg, col_reg}==14'b10101101011101)) color_data = 12'b000000001110;

		if(({row_reg, col_reg}>=14'b10101101011110) && ({row_reg, col_reg}<14'b10101110101001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==14'b10101110101001)) color_data = 12'b000000001110;
		if(({row_reg, col_reg}==14'b10101110101010)) color_data = 12'b000000001101;
		if(({row_reg, col_reg}==14'b10101110101011)) color_data = 12'b000100001101;
		if(({row_reg, col_reg}==14'b10101110101100)) color_data = 12'b000100001100;
		if(({row_reg, col_reg}==14'b10101110101101)) color_data = 12'b001000011010;
		if(({row_reg, col_reg}==14'b10101110101110)) color_data = 12'b001100101001;
		if(({row_reg, col_reg}==14'b10101110101111)) color_data = 12'b010100111000;
		if(({row_reg, col_reg}==14'b10101110110000)) color_data = 12'b010101001000;
		if(({row_reg, col_reg}==14'b10101110110001)) color_data = 12'b010101000111;
		if(({row_reg, col_reg}==14'b10101110110010)) color_data = 12'b010100110110;
		if(({row_reg, col_reg}>=14'b10101110110011) && ({row_reg, col_reg}<14'b10101110110101)) color_data = 12'b010101000111;
		if(({row_reg, col_reg}==14'b10101110110101)) color_data = 12'b010000110110;
		if(({row_reg, col_reg}==14'b10101110110110)) color_data = 12'b010100110110;
		if(({row_reg, col_reg}==14'b10101110110111)) color_data = 12'b010000110101;
		if(({row_reg, col_reg}==14'b10101110111000)) color_data = 12'b010000110100;
		if(({row_reg, col_reg}==14'b10101110111001)) color_data = 12'b101010011010;
		if(({row_reg, col_reg}==14'b10101110111010)) color_data = 12'b110010111100;
		if(({row_reg, col_reg}>=14'b10101110111011) && ({row_reg, col_reg}<14'b10101110111101)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==14'b10101110111101)) color_data = 12'b101110101001;
		if(({row_reg, col_reg}==14'b10101110111110)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==14'b10101110111111)) color_data = 12'b100001111000;
		if(({row_reg, col_reg}==14'b10101111000000)) color_data = 12'b010000100011;
		if(({row_reg, col_reg}==14'b10101111000001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=14'b10101111000010) && ({row_reg, col_reg}<14'b10101111000100)) color_data = 12'b001100010001;
		if(({row_reg, col_reg}==14'b10101111000100)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==14'b10101111000101)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==14'b10101111000110)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}>=14'b10101111000111) && ({row_reg, col_reg}<14'b10101111001001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==14'b10101111001001)) color_data = 12'b010000110011;
		if(({row_reg, col_reg}>=14'b10101111001010) && ({row_reg, col_reg}<14'b10101111001100)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}>=14'b10101111001100) && ({row_reg, col_reg}<14'b10101111001110)) color_data = 12'b010000100011;
		if(({row_reg, col_reg}>=14'b10101111001110) && ({row_reg, col_reg}<14'b10101111010000)) color_data = 12'b001100010001;
		if(({row_reg, col_reg}==14'b10101111010000)) color_data = 12'b011101010101;
		if(({row_reg, col_reg}==14'b10101111010001)) color_data = 12'b100101111000;
		if(({row_reg, col_reg}==14'b10101111010010)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==14'b10101111010011)) color_data = 12'b100101111000;
		if(({row_reg, col_reg}==14'b10101111010100)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==14'b10101111010101)) color_data = 12'b100101111000;
		if(({row_reg, col_reg}==14'b10101111010110)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==14'b10101111010111)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}>=14'b10101111011000) && ({row_reg, col_reg}<14'b10101111011010)) color_data = 12'b101110101011;
		if(({row_reg, col_reg}==14'b10101111011010)) color_data = 12'b101010011101;
		if(({row_reg, col_reg}==14'b10101111011011)) color_data = 12'b011101101101;
		if(({row_reg, col_reg}==14'b10101111011100)) color_data = 12'b001000101100;
		if(({row_reg, col_reg}==14'b10101111011101)) color_data = 12'b000000001101;

		if(({row_reg, col_reg}>=14'b10101111011110) && ({row_reg, col_reg}<14'b10110000101000)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==14'b10110000101000)) color_data = 12'b000000001110;
		if(({row_reg, col_reg}==14'b10110000101001)) color_data = 12'b000100001100;
		if(({row_reg, col_reg}==14'b10110000101010)) color_data = 12'b000100001011;
		if(({row_reg, col_reg}==14'b10110000101011)) color_data = 12'b001000011011;
		if(({row_reg, col_reg}==14'b10110000101100)) color_data = 12'b001000011010;
		if(({row_reg, col_reg}==14'b10110000101101)) color_data = 12'b010000101001;
		if(({row_reg, col_reg}==14'b10110000101110)) color_data = 12'b010100111000;
		if(({row_reg, col_reg}==14'b10110000101111)) color_data = 12'b011001000111;
		if(({row_reg, col_reg}==14'b10110000110000)) color_data = 12'b010000100110;
		if(({row_reg, col_reg}==14'b10110000110001)) color_data = 12'b010000110110;
		if(({row_reg, col_reg}==14'b10110000110010)) color_data = 12'b010000100101;
		if(({row_reg, col_reg}==14'b10110000110011)) color_data = 12'b001100100101;
		if(({row_reg, col_reg}==14'b10110000110100)) color_data = 12'b011101011000;
		if(({row_reg, col_reg}==14'b10110000110101)) color_data = 12'b110010111101;
		if(({row_reg, col_reg}==14'b10110000110110)) color_data = 12'b101110101100;
		if(({row_reg, col_reg}>=14'b10110000110111) && ({row_reg, col_reg}<14'b10110000111010)) color_data = 12'b101110101011;
		if(({row_reg, col_reg}==14'b10110000111010)) color_data = 12'b110010111011;
		if(({row_reg, col_reg}==14'b10110000111011)) color_data = 12'b101010011010;
		if(({row_reg, col_reg}==14'b10110000111100)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}>=14'b10110000111101) && ({row_reg, col_reg}<14'b10110001000000)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==14'b10110001000000)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==14'b10110001000001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=14'b10110001000010) && ({row_reg, col_reg}<14'b10110001000101)) color_data = 12'b001100010001;
		if(({row_reg, col_reg}>=14'b10110001000101) && ({row_reg, col_reg}<14'b10110001000111)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}==14'b10110001000111)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==14'b10110001001000)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}==14'b10110001001001)) color_data = 12'b010000110011;
		if(({row_reg, col_reg}==14'b10110001001010)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}>=14'b10110001001011) && ({row_reg, col_reg}<14'b10110001001101)) color_data = 12'b010000100011;
		if(({row_reg, col_reg}>=14'b10110001001101) && ({row_reg, col_reg}<14'b10110001010000)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}==14'b10110001010000)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}>=14'b10110001010001) && ({row_reg, col_reg}<14'b10110001010011)) color_data = 12'b001100010010;
		if(({row_reg, col_reg}==14'b10110001010011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==14'b10110001010100)) color_data = 12'b010000100011;
		if(({row_reg, col_reg}==14'b10110001010101)) color_data = 12'b100101111000;
		if(({row_reg, col_reg}==14'b10110001010110)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==14'b10110001010111)) color_data = 12'b100110000111;
		if(({row_reg, col_reg}>=14'b10110001011000) && ({row_reg, col_reg}<14'b10110001011010)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==14'b10110001011010)) color_data = 12'b100001111001;
		if(({row_reg, col_reg}==14'b10110001011011)) color_data = 12'b100001111011;
		if(({row_reg, col_reg}==14'b10110001011100)) color_data = 12'b010101011101;
		if(({row_reg, col_reg}==14'b10110001011101)) color_data = 12'b001000101101;
		if(({row_reg, col_reg}==14'b10110001011110)) color_data = 12'b000000001110;

		if(({row_reg, col_reg}>=14'b10110001011111) && ({row_reg, col_reg}<14'b10110010100100)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=14'b10110010100100) && ({row_reg, col_reg}<14'b10110010100111)) color_data = 12'b000000001110;
		if(({row_reg, col_reg}==14'b10110010100111)) color_data = 12'b000100001101;
		if(({row_reg, col_reg}==14'b10110010101000)) color_data = 12'b000100001011;
		if(({row_reg, col_reg}==14'b10110010101001)) color_data = 12'b001000001010;
		if(({row_reg, col_reg}==14'b10110010101010)) color_data = 12'b001100101010;
		if(({row_reg, col_reg}>=14'b10110010101011) && ({row_reg, col_reg}<14'b10110010101101)) color_data = 12'b010100111010;
		if(({row_reg, col_reg}==14'b10110010101101)) color_data = 12'b010101001001;
		if(({row_reg, col_reg}==14'b10110010101110)) color_data = 12'b011001000111;
		if(({row_reg, col_reg}==14'b10110010101111)) color_data = 12'b010101000101;
		if(({row_reg, col_reg}==14'b10110010110000)) color_data = 12'b001100100101;
		if(({row_reg, col_reg}>=14'b10110010110001) && ({row_reg, col_reg}<14'b10110010110011)) color_data = 12'b010000100101;
		if(({row_reg, col_reg}==14'b10110010110011)) color_data = 12'b001100100100;
		if(({row_reg, col_reg}==14'b10110010110100)) color_data = 12'b011001010111;
		if(({row_reg, col_reg}==14'b10110010110101)) color_data = 12'b101110101100;
		if(({row_reg, col_reg}>=14'b10110010110110) && ({row_reg, col_reg}<14'b10110010111010)) color_data = 12'b101110101011;
		if(({row_reg, col_reg}==14'b10110010111010)) color_data = 12'b110010111011;
		if(({row_reg, col_reg}==14'b10110010111011)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}>=14'b10110010111100) && ({row_reg, col_reg}<14'b10110010111110)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==14'b10110010111110)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==14'b10110010111111)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==14'b10110011000000)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}==14'b10110011000001)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=14'b10110011000010) && ({row_reg, col_reg}<14'b10110011000101)) color_data = 12'b001100010001;
		if(({row_reg, col_reg}>=14'b10110011000101) && ({row_reg, col_reg}<14'b10110011001011)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}==14'b10110011001011)) color_data = 12'b010000110011;
		if(({row_reg, col_reg}==14'b10110011001100)) color_data = 12'b010100110011;
		if(({row_reg, col_reg}==14'b10110011001101)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}>=14'b10110011001110) && ({row_reg, col_reg}<14'b10110011010000)) color_data = 12'b010100110011;
		if(({row_reg, col_reg}==14'b10110011010000)) color_data = 12'b001100010001;
		if(({row_reg, col_reg}>=14'b10110011010001) && ({row_reg, col_reg}<14'b10110011010100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==14'b10110011010100)) color_data = 12'b010000110011;
		if(({row_reg, col_reg}==14'b10110011010101)) color_data = 12'b100101111000;
		if(({row_reg, col_reg}>=14'b10110011010110) && ({row_reg, col_reg}<14'b10110011011000)) color_data = 12'b101010001000;
		if(({row_reg, col_reg}>=14'b10110011011000) && ({row_reg, col_reg}<14'b10110011011011)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==14'b10110011011011)) color_data = 12'b100110001010;
		if(({row_reg, col_reg}==14'b10110011011100)) color_data = 12'b011101111101;
		if(({row_reg, col_reg}==14'b10110011011101)) color_data = 12'b010000111101;
		if(({row_reg, col_reg}==14'b10110011011110)) color_data = 12'b000000001101;
		if(({row_reg, col_reg}==14'b10110011011111)) color_data = 12'b000000001110;

		if(({row_reg, col_reg}>=14'b10110011100000) && ({row_reg, col_reg}<14'b10110100100011)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==14'b10110100100011)) color_data = 12'b000000001110;
		if(({row_reg, col_reg}==14'b10110100100100)) color_data = 12'b000000001101;
		if(({row_reg, col_reg}==14'b10110100100101)) color_data = 12'b000100001100;
		if(({row_reg, col_reg}==14'b10110100100110)) color_data = 12'b001000011100;
		if(({row_reg, col_reg}==14'b10110100100111)) color_data = 12'b001000011010;
		if(({row_reg, col_reg}==14'b10110100101000)) color_data = 12'b001100101001;
		if(({row_reg, col_reg}==14'b10110100101001)) color_data = 12'b010000101000;
		if(({row_reg, col_reg}>=14'b10110100101010) && ({row_reg, col_reg}<14'b10110100101100)) color_data = 12'b010100111000;
		if(({row_reg, col_reg}==14'b10110100101100)) color_data = 12'b010000101000;
		if(({row_reg, col_reg}==14'b10110100101101)) color_data = 12'b010000100111;
		if(({row_reg, col_reg}==14'b10110100101110)) color_data = 12'b010000110111;
		if(({row_reg, col_reg}==14'b10110100101111)) color_data = 12'b010100110110;
		if(({row_reg, col_reg}==14'b10110100110000)) color_data = 12'b100110001010;
		if(({row_reg, col_reg}==14'b10110100110001)) color_data = 12'b101010001011;
		if(({row_reg, col_reg}==14'b10110100110010)) color_data = 12'b101010001010;
		if(({row_reg, col_reg}==14'b10110100110011)) color_data = 12'b100110001010;
		if(({row_reg, col_reg}==14'b10110100110100)) color_data = 12'b101010011010;
		if(({row_reg, col_reg}==14'b10110100110101)) color_data = 12'b110010111100;
		if(({row_reg, col_reg}>=14'b10110100110110) && ({row_reg, col_reg}<14'b10110100111000)) color_data = 12'b101110101011;
		if(({row_reg, col_reg}==14'b10110100111000)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==14'b10110100111001)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==14'b10110100111010)) color_data = 12'b100110001001;
		if(({row_reg, col_reg}>=14'b10110100111011) && ({row_reg, col_reg}<14'b10110100111101)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==14'b10110100111101)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==14'b10110100111110)) color_data = 12'b010100110011;
		if(({row_reg, col_reg}==14'b10110100111111)) color_data = 12'b010000110011;
		if(({row_reg, col_reg}==14'b10110101000000)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==14'b10110101000001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==14'b10110101000010)) color_data = 12'b001100010001;
		if(({row_reg, col_reg}>=14'b10110101000011) && ({row_reg, col_reg}<14'b10110101000101)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}==14'b10110101000101)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=14'b10110101000110) && ({row_reg, col_reg}<14'b10110101001000)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}>=14'b10110101001000) && ({row_reg, col_reg}<14'b10110101001011)) color_data = 12'b001100010001;
		if(({row_reg, col_reg}==14'b10110101001011)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}==14'b10110101001100)) color_data = 12'b010000100011;
		if(({row_reg, col_reg}>=14'b10110101001101) && ({row_reg, col_reg}<14'b10110101010000)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}==14'b10110101010000)) color_data = 12'b010000100011;
		if(({row_reg, col_reg}==14'b10110101010001)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}==14'b10110101010010)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}>=14'b10110101010011) && ({row_reg, col_reg}<14'b10110101010101)) color_data = 12'b001100010001;
		if(({row_reg, col_reg}==14'b10110101010101)) color_data = 12'b010100110011;
		if(({row_reg, col_reg}==14'b10110101010110)) color_data = 12'b010000100011;
		if(({row_reg, col_reg}==14'b10110101010111)) color_data = 12'b010000110011;
		if(({row_reg, col_reg}==14'b10110101011000)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==14'b10110101011001)) color_data = 12'b011101010101;
		if(({row_reg, col_reg}==14'b10110101011010)) color_data = 12'b100110000111;
		if(({row_reg, col_reg}==14'b10110101011011)) color_data = 12'b100110001001;
		if(({row_reg, col_reg}==14'b10110101011100)) color_data = 12'b011101101011;
		if(({row_reg, col_reg}==14'b10110101011101)) color_data = 12'b010000111100;
		if(({row_reg, col_reg}==14'b10110101011110)) color_data = 12'b000100001101;

		if(({row_reg, col_reg}>=14'b10110101011111) && ({row_reg, col_reg}<14'b10110110100001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==14'b10110110100001)) color_data = 12'b000000001110;
		if(({row_reg, col_reg}==14'b10110110100010)) color_data = 12'b000000001101;
		if(({row_reg, col_reg}==14'b10110110100011)) color_data = 12'b000100001100;
		if(({row_reg, col_reg}==14'b10110110100100)) color_data = 12'b000100001010;
		if(({row_reg, col_reg}==14'b10110110100101)) color_data = 12'b000100001001;
		if(({row_reg, col_reg}==14'b10110110100110)) color_data = 12'b001100101001;
		if(({row_reg, col_reg}==14'b10110110100111)) color_data = 12'b010000111001;
		if(({row_reg, col_reg}==14'b10110110101000)) color_data = 12'b010100111000;
		if(({row_reg, col_reg}==14'b10110110101001)) color_data = 12'b011001001000;
		if(({row_reg, col_reg}==14'b10110110101010)) color_data = 12'b010101001000;
		if(({row_reg, col_reg}==14'b10110110101011)) color_data = 12'b001100100111;
		if(({row_reg, col_reg}==14'b10110110101100)) color_data = 12'b001000010111;
		if(({row_reg, col_reg}==14'b10110110101101)) color_data = 12'b001000000111;
		if(({row_reg, col_reg}>=14'b10110110101110) && ({row_reg, col_reg}<14'b10110110110000)) color_data = 12'b001000010110;
		if(({row_reg, col_reg}==14'b10110110110000)) color_data = 12'b101110011011;
		if(({row_reg, col_reg}==14'b10110110110001)) color_data = 12'b110010101100;
		if(({row_reg, col_reg}==14'b10110110110010)) color_data = 12'b110010111100;
		if(({row_reg, col_reg}==14'b10110110110011)) color_data = 12'b110010101100;
		if(({row_reg, col_reg}==14'b10110110110100)) color_data = 12'b101110101011;
		if(({row_reg, col_reg}==14'b10110110110101)) color_data = 12'b110010111011;
		if(({row_reg, col_reg}>=14'b10110110110110) && ({row_reg, col_reg}<14'b10110110111000)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==14'b10110110111000)) color_data = 12'b110010111011;
		if(({row_reg, col_reg}==14'b10110110111001)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==14'b10110110111010)) color_data = 12'b100001111000;
		if(({row_reg, col_reg}==14'b10110110111011)) color_data = 12'b100101111000;
		if(({row_reg, col_reg}==14'b10110110111100)) color_data = 12'b100110001001;
		if(({row_reg, col_reg}==14'b10110110111101)) color_data = 12'b100001100110;
		if(({row_reg, col_reg}==14'b10110110111110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==14'b10110110111111)) color_data = 12'b001000000000;
		if(({row_reg, col_reg}==14'b10110111000000)) color_data = 12'b001100010001;
		if(({row_reg, col_reg}==14'b10110111000001)) color_data = 12'b001000000000;
		if(({row_reg, col_reg}==14'b10110111000010)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}==14'b10110111000011)) color_data = 12'b010100110011;
		if(({row_reg, col_reg}==14'b10110111000100)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}==14'b10110111000101)) color_data = 12'b010100100010;
		if(({row_reg, col_reg}==14'b10110111000110)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}>=14'b10110111000111) && ({row_reg, col_reg}<14'b10110111001011)) color_data = 12'b001100010001;
		if(({row_reg, col_reg}==14'b10110111001011)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}>=14'b10110111001100) && ({row_reg, col_reg}<14'b10110111001110)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}==14'b10110111001110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=14'b10110111001111) && ({row_reg, col_reg}<14'b10110111010011)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}>=14'b10110111010011) && ({row_reg, col_reg}<14'b10110111010110)) color_data = 12'b001100010001;
		if(({row_reg, col_reg}==14'b10110111010110)) color_data = 12'b001000000000;
		if(({row_reg, col_reg}==14'b10110111010111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==14'b10110111011000)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==14'b10110111011001)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==14'b10110111011010)) color_data = 12'b101010001000;
		if(({row_reg, col_reg}==14'b10110111011011)) color_data = 12'b101010011010;
		if(({row_reg, col_reg}==14'b10110111011100)) color_data = 12'b100001111011;
		if(({row_reg, col_reg}==14'b10110111011101)) color_data = 12'b010000111011;
		if(({row_reg, col_reg}==14'b10110111011110)) color_data = 12'b000100011101;
		if(({row_reg, col_reg}==14'b10110111011111)) color_data = 12'b000000001110;

		if(({row_reg, col_reg}>=14'b10110111100000) && ({row_reg, col_reg}<14'b10111000011110)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=14'b10111000011110) && ({row_reg, col_reg}<14'b10111000100000)) color_data = 12'b000000001110;
		if(({row_reg, col_reg}==14'b10111000100000)) color_data = 12'b000000001101;
		if(({row_reg, col_reg}==14'b10111000100001)) color_data = 12'b000100001100;
		if(({row_reg, col_reg}==14'b10111000100010)) color_data = 12'b000100001011;
		if(({row_reg, col_reg}==14'b10111000100011)) color_data = 12'b001000011010;
		if(({row_reg, col_reg}==14'b10111000100100)) color_data = 12'b001100101001;
		if(({row_reg, col_reg}==14'b10111000100101)) color_data = 12'b010000101001;
		if(({row_reg, col_reg}==14'b10111000100110)) color_data = 12'b010101001001;
		if(({row_reg, col_reg}==14'b10111000100111)) color_data = 12'b010101001000;
		if(({row_reg, col_reg}>=14'b10111000101000) && ({row_reg, col_reg}<14'b10111000101010)) color_data = 12'b010000110111;
		if(({row_reg, col_reg}==14'b10111000101010)) color_data = 12'b001100100111;
		if(({row_reg, col_reg}==14'b10111000101011)) color_data = 12'b001000011000;
		if(({row_reg, col_reg}>=14'b10111000101100) && ({row_reg, col_reg}<14'b10111000101110)) color_data = 12'b000100011001;
		if(({row_reg, col_reg}==14'b10111000101110)) color_data = 12'b001000011001;
		if(({row_reg, col_reg}==14'b10111000101111)) color_data = 12'b001100101001;
		if(({row_reg, col_reg}==14'b10111000110000)) color_data = 12'b101110101011;
		if(({row_reg, col_reg}>=14'b10111000110001) && ({row_reg, col_reg}<14'b10111000110011)) color_data = 12'b110010101011;
		if(({row_reg, col_reg}==14'b10111000110011)) color_data = 12'b110010111011;
		if(({row_reg, col_reg}==14'b10111000110100)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==14'b10111000110101)) color_data = 12'b101110101011;
		if(({row_reg, col_reg}==14'b10111000110110)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}>=14'b10111000110111) && ({row_reg, col_reg}<14'b10111000111001)) color_data = 12'b110010101011;
		if(({row_reg, col_reg}==14'b10111000111001)) color_data = 12'b101010001001;
		if(({row_reg, col_reg}>=14'b10111000111010) && ({row_reg, col_reg}<14'b10111000111100)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==14'b10111000111100)) color_data = 12'b101010001001;
		if(({row_reg, col_reg}==14'b10111000111101)) color_data = 12'b100001100111;
		if(({row_reg, col_reg}>=14'b10111000111110) && ({row_reg, col_reg}<14'b10111001000010)) color_data = 12'b001100010001;
		if(({row_reg, col_reg}>=14'b10111001000010) && ({row_reg, col_reg}<14'b10111001000101)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}==14'b10111001000101)) color_data = 12'b010100100010;
		if(({row_reg, col_reg}==14'b10111001000110)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}>=14'b10111001000111) && ({row_reg, col_reg}<14'b10111001001100)) color_data = 12'b001100010001;
		if(({row_reg, col_reg}==14'b10111001001100)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}>=14'b10111001001101) && ({row_reg, col_reg}<14'b10111001010001)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}==14'b10111001010001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=14'b10111001010010) && ({row_reg, col_reg}<14'b10111001010100)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}==14'b10111001010100)) color_data = 12'b001100010001;
		if(({row_reg, col_reg}==14'b10111001010101)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}==14'b10111001010110)) color_data = 12'b001100010010;
		if(({row_reg, col_reg}==14'b10111001010111)) color_data = 12'b010000100011;
		if(({row_reg, col_reg}==14'b10111001011000)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==14'b10111001011001)) color_data = 12'b010101000100;
		if(({row_reg, col_reg}==14'b10111001011010)) color_data = 12'b011001010100;
		if(({row_reg, col_reg}==14'b10111001011011)) color_data = 12'b011001010101;
		if(({row_reg, col_reg}==14'b10111001011100)) color_data = 12'b010101000111;
		if(({row_reg, col_reg}==14'b10111001011101)) color_data = 12'b001100101001;
		if(({row_reg, col_reg}==14'b10111001011110)) color_data = 12'b000100001011;
		if(({row_reg, col_reg}==14'b10111001011111)) color_data = 12'b000000001101;

		if(({row_reg, col_reg}>=14'b10111001100000) && ({row_reg, col_reg}<14'b10111010011100)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==14'b10111010011100)) color_data = 12'b000000001110;
		if(({row_reg, col_reg}>=14'b10111010011101) && ({row_reg, col_reg}<14'b10111010100000)) color_data = 12'b000000001101;
		if(({row_reg, col_reg}==14'b10111010100000)) color_data = 12'b000000001001;
		if(({row_reg, col_reg}==14'b10111010100001)) color_data = 12'b001000011010;
		if(({row_reg, col_reg}==14'b10111010100010)) color_data = 12'b001000011001;
		if(({row_reg, col_reg}==14'b10111010100011)) color_data = 12'b001100101000;
		if(({row_reg, col_reg}==14'b10111010100100)) color_data = 12'b010000111001;
		if(({row_reg, col_reg}==14'b10111010100101)) color_data = 12'b010101001001;
		if(({row_reg, col_reg}==14'b10111010100110)) color_data = 12'b010100111001;
		if(({row_reg, col_reg}==14'b10111010100111)) color_data = 12'b001100100111;
		if(({row_reg, col_reg}==14'b10111010101000)) color_data = 12'b001000010111;
		if(({row_reg, col_reg}==14'b10111010101001)) color_data = 12'b000100011000;
		if(({row_reg, col_reg}==14'b10111010101010)) color_data = 12'b000000001000;
		if(({row_reg, col_reg}==14'b10111010101011)) color_data = 12'b000000001010;
		if(({row_reg, col_reg}==14'b10111010101100)) color_data = 12'b000100001100;
		if(({row_reg, col_reg}==14'b10111010101101)) color_data = 12'b000100001011;
		if(({row_reg, col_reg}==14'b10111010101110)) color_data = 12'b001100101011;
		if(({row_reg, col_reg}==14'b10111010101111)) color_data = 12'b011001011101;
		if(({row_reg, col_reg}>=14'b10111010110000) && ({row_reg, col_reg}<14'b10111010110010)) color_data = 12'b101110101011;
		if(({row_reg, col_reg}==14'b10111010110010)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==14'b10111010110011)) color_data = 12'b110010111011;
		if(({row_reg, col_reg}==14'b10111010110100)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==14'b10111010110101)) color_data = 12'b110010101011;
		if(({row_reg, col_reg}>=14'b10111010110110) && ({row_reg, col_reg}<14'b10111010111000)) color_data = 12'b110010111011;
		if(({row_reg, col_reg}==14'b10111010111000)) color_data = 12'b101110101011;
		if(({row_reg, col_reg}==14'b10111010111001)) color_data = 12'b101010001001;
		if(({row_reg, col_reg}>=14'b10111010111010) && ({row_reg, col_reg}<14'b10111010111100)) color_data = 12'b100101111000;
		if(({row_reg, col_reg}==14'b10111010111100)) color_data = 12'b100110001001;
		if(({row_reg, col_reg}==14'b10111010111101)) color_data = 12'b100001100111;
		if(({row_reg, col_reg}>=14'b10111010111110) && ({row_reg, col_reg}<14'b10111011000010)) color_data = 12'b001100010001;
		if(({row_reg, col_reg}>=14'b10111011000010) && ({row_reg, col_reg}<14'b10111011000101)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}==14'b10111011000101)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==14'b10111011000110)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}==14'b10111011000111)) color_data = 12'b001100010001;
		if(({row_reg, col_reg}==14'b10111011001000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=14'b10111011001001) && ({row_reg, col_reg}<14'b10111011001011)) color_data = 12'b001100010001;
		if(({row_reg, col_reg}==14'b10111011001011)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=14'b10111011001100) && ({row_reg, col_reg}<14'b10111011001110)) color_data = 12'b001100010001;
		if(({row_reg, col_reg}>=14'b10111011001110) && ({row_reg, col_reg}<14'b10111011010101)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}==14'b10111011010101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==14'b10111011010110)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}>=14'b10111011010111) && ({row_reg, col_reg}<14'b10111011011001)) color_data = 12'b010000110011;
		if(({row_reg, col_reg}==14'b10111011011001)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}>=14'b10111011011010) && ({row_reg, col_reg}<14'b10111011011100)) color_data = 12'b001000000000;
		if(({row_reg, col_reg}==14'b10111011011100)) color_data = 12'b001000000010;
		if(({row_reg, col_reg}==14'b10111011011101)) color_data = 12'b000100000101;
		if(({row_reg, col_reg}==14'b10111011011110)) color_data = 12'b000000001001;
		if(({row_reg, col_reg}==14'b10111011011111)) color_data = 12'b000100001100;

		if(({row_reg, col_reg}>=14'b10111011100000) && ({row_reg, col_reg}<14'b10111100011010)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==14'b10111100011010)) color_data = 12'b000000001110;
		if(({row_reg, col_reg}==14'b10111100011011)) color_data = 12'b000000001101;
		if(({row_reg, col_reg}>=14'b10111100011100) && ({row_reg, col_reg}<14'b10111100011110)) color_data = 12'b000000001100;
		if(({row_reg, col_reg}==14'b10111100011110)) color_data = 12'b000100001011;
		if(({row_reg, col_reg}==14'b10111100011111)) color_data = 12'b000100011011;
		if(({row_reg, col_reg}==14'b10111100100000)) color_data = 12'b001100011000;
		if(({row_reg, col_reg}>=14'b10111100100001) && ({row_reg, col_reg}<14'b10111100100011)) color_data = 12'b010000111001;
		if(({row_reg, col_reg}==14'b10111100100011)) color_data = 12'b010100111000;
		if(({row_reg, col_reg}==14'b10111100100100)) color_data = 12'b010101001001;
		if(({row_reg, col_reg}==14'b10111100100101)) color_data = 12'b010100111001;
		if(({row_reg, col_reg}==14'b10111100100110)) color_data = 12'b001100101001;
		if(({row_reg, col_reg}==14'b10111100100111)) color_data = 12'b001000011001;
		if(({row_reg, col_reg}==14'b10111100101000)) color_data = 12'b000100001001;
		if(({row_reg, col_reg}==14'b10111100101001)) color_data = 12'b000000001010;
		if(({row_reg, col_reg}==14'b10111100101010)) color_data = 12'b000000001100;
		if(({row_reg, col_reg}==14'b10111100101011)) color_data = 12'b000000001110;
		if(({row_reg, col_reg}==14'b10111100101100)) color_data = 12'b000000001101;
		if(({row_reg, col_reg}==14'b10111100101101)) color_data = 12'b000000001011;
		if(({row_reg, col_reg}==14'b10111100101110)) color_data = 12'b001100101011;
		if(({row_reg, col_reg}==14'b10111100101111)) color_data = 12'b011101101101;
		if(({row_reg, col_reg}>=14'b10111100110000) && ({row_reg, col_reg}<14'b10111100110010)) color_data = 12'b101110101011;
		if(({row_reg, col_reg}==14'b10111100110010)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==14'b10111100110011)) color_data = 12'b110010111011;
		if(({row_reg, col_reg}==14'b10111100110100)) color_data = 12'b110010101010;
		if(({row_reg, col_reg}==14'b10111100110101)) color_data = 12'b110010111011;
		if(({row_reg, col_reg}==14'b10111100110110)) color_data = 12'b110010101011;
		if(({row_reg, col_reg}==14'b10111100110111)) color_data = 12'b101110011010;
		if(({row_reg, col_reg}==14'b10111100111000)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==14'b10111100111001)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}>=14'b10111100111010) && ({row_reg, col_reg}<14'b10111100111100)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==14'b10111100111100)) color_data = 12'b101010001001;
		if(({row_reg, col_reg}==14'b10111100111101)) color_data = 12'b100001100111;
		if(({row_reg, col_reg}==14'b10111100111110)) color_data = 12'b001100010001;
		if(({row_reg, col_reg}==14'b10111100111111)) color_data = 12'b001100010000;
		if(({row_reg, col_reg}>=14'b10111101000000) && ({row_reg, col_reg}<14'b10111101000010)) color_data = 12'b001100010001;
		if(({row_reg, col_reg}>=14'b10111101000010) && ({row_reg, col_reg}<14'b10111101000100)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}==14'b10111101000100)) color_data = 12'b010100100010;
		if(({row_reg, col_reg}>=14'b10111101000101) && ({row_reg, col_reg}<14'b10111101001000)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}==14'b10111101001000)) color_data = 12'b001100010001;
		if(({row_reg, col_reg}==14'b10111101001001)) color_data = 12'b001100010010;
		if(({row_reg, col_reg}>=14'b10111101001010) && ({row_reg, col_reg}<14'b10111101001100)) color_data = 12'b001100010001;
		if(({row_reg, col_reg}==14'b10111101001100)) color_data = 12'b001100010010;
		if(({row_reg, col_reg}==14'b10111101001101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=14'b10111101001110) && ({row_reg, col_reg}<14'b10111101010001)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}==14'b10111101010001)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}==14'b10111101010010)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}==14'b10111101010011)) color_data = 12'b010100110011;
		if(({row_reg, col_reg}==14'b10111101010100)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}==14'b10111101010101)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==14'b10111101010110)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}==14'b10111101010111)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==14'b10111101011000)) color_data = 12'b010000100011;
		if(({row_reg, col_reg}==14'b10111101011001)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}>=14'b10111101011010) && ({row_reg, col_reg}<14'b10111101011100)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==14'b10111101011100)) color_data = 12'b001100010010;
		if(({row_reg, col_reg}==14'b10111101011101)) color_data = 12'b000100000100;
		if(({row_reg, col_reg}==14'b10111101011110)) color_data = 12'b000100001000;
		if(({row_reg, col_reg}==14'b10111101011111)) color_data = 12'b000100001011;

		if(({row_reg, col_reg}>=14'b10111101100000) && ({row_reg, col_reg}<14'b10111110011010)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==14'b10111110011010)) color_data = 12'b000000001110;
		if(({row_reg, col_reg}==14'b10111110011011)) color_data = 12'b000000001101;
		if(({row_reg, col_reg}==14'b10111110011100)) color_data = 12'b000000001100;
		if(({row_reg, col_reg}==14'b10111110011101)) color_data = 12'b000100001011;
		if(({row_reg, col_reg}==14'b10111110011110)) color_data = 12'b000100011010;
		if(({row_reg, col_reg}==14'b10111110011111)) color_data = 12'b001000011010;
		if(({row_reg, col_reg}==14'b10111110100000)) color_data = 12'b010000110111;
		if(({row_reg, col_reg}==14'b10111110100001)) color_data = 12'b010101001001;
		if(({row_reg, col_reg}==14'b10111110100010)) color_data = 12'b010000110111;
		if(({row_reg, col_reg}==14'b10111110100011)) color_data = 12'b010000100111;
		if(({row_reg, col_reg}==14'b10111110100100)) color_data = 12'b001100100111;
		if(({row_reg, col_reg}==14'b10111110100101)) color_data = 12'b001000010111;
		if(({row_reg, col_reg}==14'b10111110100110)) color_data = 12'b000100001000;
		if(({row_reg, col_reg}==14'b10111110100111)) color_data = 12'b000100001010;
		if(({row_reg, col_reg}==14'b10111110101000)) color_data = 12'b000000001100;
		if(({row_reg, col_reg}==14'b10111110101001)) color_data = 12'b000000001101;
		if(({row_reg, col_reg}>=14'b10111110101010) && ({row_reg, col_reg}<14'b10111110101101)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==14'b10111110101101)) color_data = 12'b000100001100;
		if(({row_reg, col_reg}==14'b10111110101110)) color_data = 12'b010001001100;
		if(({row_reg, col_reg}==14'b10111110101111)) color_data = 12'b100110001101;
		if(({row_reg, col_reg}==14'b10111110110000)) color_data = 12'b110010101100;
		if(({row_reg, col_reg}==14'b10111110110001)) color_data = 12'b110010111011;
		if(({row_reg, col_reg}==14'b10111110110010)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==14'b10111110110011)) color_data = 12'b110010111011;
		if(({row_reg, col_reg}==14'b10111110110100)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==14'b10111110110101)) color_data = 12'b110010101011;
		if(({row_reg, col_reg}==14'b10111110110110)) color_data = 12'b101110101011;
		if(({row_reg, col_reg}==14'b10111110110111)) color_data = 12'b100110001001;
		if(({row_reg, col_reg}==14'b10111110111000)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==14'b10111110111001)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}>=14'b10111110111010) && ({row_reg, col_reg}<14'b10111110111100)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==14'b10111110111100)) color_data = 12'b100110001001;
		if(({row_reg, col_reg}==14'b10111110111101)) color_data = 12'b100001100111;
		if(({row_reg, col_reg}==14'b10111110111110)) color_data = 12'b001100010001;
		if(({row_reg, col_reg}==14'b10111110111111)) color_data = 12'b001100010000;
		if(({row_reg, col_reg}>=14'b10111111000000) && ({row_reg, col_reg}<14'b10111111000101)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}>=14'b10111111000101) && ({row_reg, col_reg}<14'b10111111000111)) color_data = 12'b001100010001;
		if(({row_reg, col_reg}==14'b10111111000111)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}==14'b10111111001000)) color_data = 12'b010000100011;
		if(({row_reg, col_reg}==14'b10111111001001)) color_data = 12'b001100010010;
		if(({row_reg, col_reg}==14'b10111111001010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==14'b10111111001011)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}>=14'b10111111001100) && ({row_reg, col_reg}<14'b10111111001110)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}>=14'b10111111001110) && ({row_reg, col_reg}<14'b10111111010000)) color_data = 12'b001100010001;
		if(({row_reg, col_reg}==14'b10111111010000)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==14'b10111111010001)) color_data = 12'b010100100010;
		if(({row_reg, col_reg}==14'b10111111010010)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}==14'b10111111010011)) color_data = 12'b010100100011;
		if(({row_reg, col_reg}>=14'b10111111010100) && ({row_reg, col_reg}<14'b10111111010110)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}==14'b10111111010110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==14'b10111111010111)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}==14'b10111111011000)) color_data = 12'b010000100011;
		if(({row_reg, col_reg}>=14'b10111111011001) && ({row_reg, col_reg}<14'b10111111011011)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}==14'b10111111011011)) color_data = 12'b010000110001;
		if(({row_reg, col_reg}==14'b10111111011100)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}==14'b10111111011101)) color_data = 12'b001100100100;
		if(({row_reg, col_reg}==14'b10111111011110)) color_data = 12'b000100000111;
		if(({row_reg, col_reg}==14'b10111111011111)) color_data = 12'b000000001000;

		if(({row_reg, col_reg}>=14'b10111111100000) && ({row_reg, col_reg}<14'b11000000011001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==14'b11000000011001)) color_data = 12'b000000001110;
		if(({row_reg, col_reg}==14'b11000000011010)) color_data = 12'b000100011100;
		if(({row_reg, col_reg}==14'b11000000011011)) color_data = 12'b000100001001;
		if(({row_reg, col_reg}==14'b11000000011100)) color_data = 12'b001100011000;
		if(({row_reg, col_reg}==14'b11000000011101)) color_data = 12'b010100111001;
		if(({row_reg, col_reg}==14'b11000000011110)) color_data = 12'b010101001000;
		if(({row_reg, col_reg}==14'b11000000011111)) color_data = 12'b011001000111;
		if(({row_reg, col_reg}==14'b11000000100000)) color_data = 12'b010101001000;
		if(({row_reg, col_reg}==14'b11000000100001)) color_data = 12'b010000111000;
		if(({row_reg, col_reg}==14'b11000000100010)) color_data = 12'b001000011000;
		if(({row_reg, col_reg}==14'b11000000100011)) color_data = 12'b000100001001;
		if(({row_reg, col_reg}==14'b11000000100100)) color_data = 12'b000000001010;
		if(({row_reg, col_reg}==14'b11000000100101)) color_data = 12'b000000001011;
		if(({row_reg, col_reg}==14'b11000000100110)) color_data = 12'b000000001100;
		if(({row_reg, col_reg}==14'b11000000100111)) color_data = 12'b000000001101;
		if(({row_reg, col_reg}>=14'b11000000101000) && ({row_reg, col_reg}<14'b11000000101010)) color_data = 12'b000000001110;
		if(({row_reg, col_reg}>=14'b11000000101010) && ({row_reg, col_reg}<14'b11000000101100)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==14'b11000000101100)) color_data = 12'b000000001110;
		if(({row_reg, col_reg}==14'b11000000101101)) color_data = 12'b001000011100;
		if(({row_reg, col_reg}==14'b11000000101110)) color_data = 12'b011001011100;
		if(({row_reg, col_reg}==14'b11000000101111)) color_data = 12'b101010011100;
		if(({row_reg, col_reg}==14'b11000000110000)) color_data = 12'b110010111011;
		if(({row_reg, col_reg}==14'b11000000110001)) color_data = 12'b101110101011;
		if(({row_reg, col_reg}>=14'b11000000110010) && ({row_reg, col_reg}<14'b11000000110101)) color_data = 12'b110010101011;
		if(({row_reg, col_reg}>=14'b11000000110101) && ({row_reg, col_reg}<14'b11000000110111)) color_data = 12'b101110101011;
		if(({row_reg, col_reg}>=14'b11000000110111) && ({row_reg, col_reg}<14'b11000000111011)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==14'b11000000111011)) color_data = 12'b100101111000;
		if(({row_reg, col_reg}==14'b11000000111100)) color_data = 12'b101010001000;
		if(({row_reg, col_reg}==14'b11000000111101)) color_data = 12'b100001100110;
		if(({row_reg, col_reg}>=14'b11000000111110) && ({row_reg, col_reg}<14'b11000001000000)) color_data = 12'b001100010001;
		if(({row_reg, col_reg}==14'b11000001000000)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}>=14'b11000001000001) && ({row_reg, col_reg}<14'b11000001000011)) color_data = 12'b010000100011;
		if(({row_reg, col_reg}>=14'b11000001000011) && ({row_reg, col_reg}<14'b11000001000101)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}>=14'b11000001000101) && ({row_reg, col_reg}<14'b11000001000111)) color_data = 12'b001100010001;
		if(({row_reg, col_reg}==14'b11000001000111)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}==14'b11000001001000)) color_data = 12'b010000110011;
		if(({row_reg, col_reg}>=14'b11000001001001) && ({row_reg, col_reg}<14'b11000001001100)) color_data = 12'b001100010001;
		if(({row_reg, col_reg}>=14'b11000001001100) && ({row_reg, col_reg}<14'b11000001001110)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}>=14'b11000001001110) && ({row_reg, col_reg}<14'b11000001010000)) color_data = 12'b001100010001;
		if(({row_reg, col_reg}>=14'b11000001010000) && ({row_reg, col_reg}<14'b11000001010010)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}==14'b11000001010010)) color_data = 12'b010000100011;
		if(({row_reg, col_reg}==14'b11000001010011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=14'b11000001010100) && ({row_reg, col_reg}<14'b11000001010111)) color_data = 12'b010100100010;
		if(({row_reg, col_reg}>=14'b11000001010111) && ({row_reg, col_reg}<14'b11000001011101)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}==14'b11000001011101)) color_data = 12'b010000100011;
		if(({row_reg, col_reg}==14'b11000001011110)) color_data = 12'b001100100100;
		if(({row_reg, col_reg}==14'b11000001011111)) color_data = 12'b000100000100;
		if(({row_reg, col_reg}==14'b11000001100000)) color_data = 12'b000000001100;
		if(({row_reg, col_reg}==14'b11000001100001)) color_data = 12'b000000001101;

		if(({row_reg, col_reg}>=14'b11000001100010) && ({row_reg, col_reg}<14'b11000010011000)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==14'b11000010011000)) color_data = 12'b000000001110;
		if(({row_reg, col_reg}==14'b11000010011001)) color_data = 12'b000000001011;
		if(({row_reg, col_reg}==14'b11000010011010)) color_data = 12'b001000011010;
		if(({row_reg, col_reg}==14'b11000010011011)) color_data = 12'b001100101010;
		if(({row_reg, col_reg}==14'b11000010011100)) color_data = 12'b010000111001;
		if(({row_reg, col_reg}==14'b11000010011101)) color_data = 12'b010100111001;
		if(({row_reg, col_reg}>=14'b11000010011110) && ({row_reg, col_reg}<14'b11000010100000)) color_data = 12'b010000101000;
		if(({row_reg, col_reg}==14'b11000010100000)) color_data = 12'b001100101000;
		if(({row_reg, col_reg}==14'b11000010100001)) color_data = 12'b001000011001;
		if(({row_reg, col_reg}==14'b11000010100010)) color_data = 12'b000100011001;
		if(({row_reg, col_reg}==14'b11000010100011)) color_data = 12'b000000001010;
		if(({row_reg, col_reg}==14'b11000010100100)) color_data = 12'b000000001100;
		if(({row_reg, col_reg}>=14'b11000010100101) && ({row_reg, col_reg}<14'b11000010100111)) color_data = 12'b000000001101;
		if(({row_reg, col_reg}>=14'b11000010100111) && ({row_reg, col_reg}<14'b11000010101010)) color_data = 12'b000000001110;
		if(({row_reg, col_reg}>=14'b11000010101010) && ({row_reg, col_reg}<14'b11000010101100)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==14'b11000010101100)) color_data = 12'b000000001110;
		if(({row_reg, col_reg}==14'b11000010101101)) color_data = 12'b001000101100;
		if(({row_reg, col_reg}==14'b11000010101110)) color_data = 12'b011101101101;
		if(({row_reg, col_reg}==14'b11000010101111)) color_data = 12'b101110101101;
		if(({row_reg, col_reg}>=14'b11000010110000) && ({row_reg, col_reg}<14'b11000010110010)) color_data = 12'b101110101011;
		if(({row_reg, col_reg}==14'b11000010110010)) color_data = 12'b110010111011;
		if(({row_reg, col_reg}>=14'b11000010110011) && ({row_reg, col_reg}<14'b11000010110111)) color_data = 12'b101110101011;
		if(({row_reg, col_reg}==14'b11000010110111)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==14'b11000010111000)) color_data = 12'b100101111000;
		if(({row_reg, col_reg}>=14'b11000010111001) && ({row_reg, col_reg}<14'b11000010111011)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==14'b11000010111011)) color_data = 12'b011001000101;
		if(({row_reg, col_reg}==14'b11000010111100)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}==14'b11000010111101)) color_data = 12'b010000100011;
		if(({row_reg, col_reg}==14'b11000010111110)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}==14'b11000010111111)) color_data = 12'b010000100011;
		if(({row_reg, col_reg}>=14'b11000011000000) && ({row_reg, col_reg}<14'b11000011000011)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}>=14'b11000011000011) && ({row_reg, col_reg}<14'b11000011001000)) color_data = 12'b001100010001;
		if(({row_reg, col_reg}==14'b11000011001000)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}>=14'b11000011001001) && ({row_reg, col_reg}<14'b11000011001100)) color_data = 12'b001100010001;
		if(({row_reg, col_reg}>=14'b11000011001100) && ({row_reg, col_reg}<14'b11000011001110)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}>=14'b11000011001110) && ({row_reg, col_reg}<14'b11000011010101)) color_data = 12'b001100010001;
		if(({row_reg, col_reg}>=14'b11000011010101) && ({row_reg, col_reg}<14'b11000011011000)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}>=14'b11000011011000) && ({row_reg, col_reg}<14'b11000011011010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=14'b11000011011010) && ({row_reg, col_reg}<14'b11000011011101)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}==14'b11000011011101)) color_data = 12'b010000110011;
		if(({row_reg, col_reg}==14'b11000011011110)) color_data = 12'b010000100101;
		if(({row_reg, col_reg}==14'b11000011011111)) color_data = 12'b000100000100;
		if(({row_reg, col_reg}==14'b11000011100000)) color_data = 12'b000000001100;
		if(({row_reg, col_reg}==14'b11000011100001)) color_data = 12'b000000001101;

		if(({row_reg, col_reg}>=14'b11000011100010) && ({row_reg, col_reg}<14'b11000100010110)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==14'b11000100010110)) color_data = 12'b000000001110;
		if(({row_reg, col_reg}==14'b11000100010111)) color_data = 12'b000000001101;
		if(({row_reg, col_reg}==14'b11000100011000)) color_data = 12'b000100001100;
		if(({row_reg, col_reg}==14'b11000100011001)) color_data = 12'b000100001001;
		if(({row_reg, col_reg}==14'b11000100011010)) color_data = 12'b001100101001;
		if(({row_reg, col_reg}>=14'b11000100011011) && ({row_reg, col_reg}<14'b11000100011101)) color_data = 12'b010101001001;
		if(({row_reg, col_reg}==14'b11000100011101)) color_data = 12'b010000101001;
		if(({row_reg, col_reg}==14'b11000100011110)) color_data = 12'b001000001000;
		if(({row_reg, col_reg}==14'b11000100011111)) color_data = 12'b000100001000;
		if(({row_reg, col_reg}==14'b11000100100000)) color_data = 12'b000100001001;
		if(({row_reg, col_reg}==14'b11000100100001)) color_data = 12'b000000001010;
		if(({row_reg, col_reg}==14'b11000100100010)) color_data = 12'b000000001100;
		if(({row_reg, col_reg}==14'b11000100100011)) color_data = 12'b000000001101;
		if(({row_reg, col_reg}>=14'b11000100100100) && ({row_reg, col_reg}<14'b11000100100111)) color_data = 12'b000000001110;
		if(({row_reg, col_reg}>=14'b11000100100111) && ({row_reg, col_reg}<14'b11000100101100)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==14'b11000100101100)) color_data = 12'b000000001101;
		if(({row_reg, col_reg}==14'b11000100101101)) color_data = 12'b001100111101;
		if(({row_reg, col_reg}==14'b11000100101110)) color_data = 12'b100001111101;
		if(({row_reg, col_reg}==14'b11000100101111)) color_data = 12'b101110101101;
		if(({row_reg, col_reg}==14'b11000100110000)) color_data = 12'b110010101011;
		if(({row_reg, col_reg}>=14'b11000100110001) && ({row_reg, col_reg}<14'b11000100110100)) color_data = 12'b101110101011;
		if(({row_reg, col_reg}==14'b11000100110100)) color_data = 12'b110010111011;
		if(({row_reg, col_reg}>=14'b11000100110101) && ({row_reg, col_reg}<14'b11000100110111)) color_data = 12'b101110101011;
		if(({row_reg, col_reg}>=14'b11000100110111) && ({row_reg, col_reg}<14'b11000100111010)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==14'b11000100111010)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==14'b11000100111011)) color_data = 12'b011001010101;
		if(({row_reg, col_reg}==14'b11000100111100)) color_data = 12'b001000000000;
		if(({row_reg, col_reg}==14'b11000100111101)) color_data = 12'b001100010001;
		if(({row_reg, col_reg}==14'b11000100111110)) color_data = 12'b010000100011;
		if(({row_reg, col_reg}==14'b11000100111111)) color_data = 12'b010100110011;
		if(({row_reg, col_reg}>=14'b11000101000000) && ({row_reg, col_reg}<14'b11000101000010)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}==14'b11000101000010)) color_data = 12'b001100010010;
		if(({row_reg, col_reg}>=14'b11000101000011) && ({row_reg, col_reg}<14'b11000101001011)) color_data = 12'b001100010001;
		if(({row_reg, col_reg}==14'b11000101001011)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}>=14'b11000101001100) && ({row_reg, col_reg}<14'b11000101001110)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}>=14'b11000101001110) && ({row_reg, col_reg}<14'b11000101010000)) color_data = 12'b001100010001;
		if(({row_reg, col_reg}==14'b11000101010000)) color_data = 12'b001100010000;
		if(({row_reg, col_reg}>=14'b11000101010001) && ({row_reg, col_reg}<14'b11000101010101)) color_data = 12'b001100010001;
		if(({row_reg, col_reg}==14'b11000101010101)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}==14'b11000101010110)) color_data = 12'b010100100011;
		if(({row_reg, col_reg}==14'b11000101010111)) color_data = 12'b010000100011;
		if(({row_reg, col_reg}==14'b11000101011000)) color_data = 12'b010000110011;
		if(({row_reg, col_reg}>=14'b11000101011001) && ({row_reg, col_reg}<14'b11000101011101)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}==14'b11000101011101)) color_data = 12'b010000110011;
		if(({row_reg, col_reg}==14'b11000101011110)) color_data = 12'b010000100100;
		if(({row_reg, col_reg}==14'b11000101011111)) color_data = 12'b000100000100;
		if(({row_reg, col_reg}==14'b11000101100000)) color_data = 12'b000000001100;
		if(({row_reg, col_reg}==14'b11000101100001)) color_data = 12'b000000001101;

		if(({row_reg, col_reg}>=14'b11000101100010) && ({row_reg, col_reg}<14'b11000110010100)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==14'b11000110010100)) color_data = 12'b000000001110;
		if(({row_reg, col_reg}==14'b11000110010101)) color_data = 12'b000000001101;
		if(({row_reg, col_reg}==14'b11000110010110)) color_data = 12'b000100001100;
		if(({row_reg, col_reg}==14'b11000110010111)) color_data = 12'b000100001011;
		if(({row_reg, col_reg}==14'b11000110011000)) color_data = 12'b001000011001;
		if(({row_reg, col_reg}==14'b11000110011001)) color_data = 12'b001100101000;
		if(({row_reg, col_reg}==14'b11000110011010)) color_data = 12'b010100111000;
		if(({row_reg, col_reg}==14'b11000110011011)) color_data = 12'b010000111000;
		if(({row_reg, col_reg}==14'b11000110011100)) color_data = 12'b001100101000;
		if(({row_reg, col_reg}==14'b11000110011101)) color_data = 12'b001000011001;
		if(({row_reg, col_reg}==14'b11000110011110)) color_data = 12'b000100001010;
		if(({row_reg, col_reg}==14'b11000110011111)) color_data = 12'b000000001010;
		if(({row_reg, col_reg}==14'b11000110100000)) color_data = 12'b000000001100;
		if(({row_reg, col_reg}==14'b11000110100001)) color_data = 12'b000000001101;
		if(({row_reg, col_reg}==14'b11000110100010)) color_data = 12'b000000001110;
		if(({row_reg, col_reg}>=14'b11000110100011) && ({row_reg, col_reg}<14'b11000110101011)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==14'b11000110101011)) color_data = 12'b000000001110;
		if(({row_reg, col_reg}==14'b11000110101100)) color_data = 12'b000100001101;
		if(({row_reg, col_reg}==14'b11000110101101)) color_data = 12'b010101001101;
		if(({row_reg, col_reg}==14'b11000110101110)) color_data = 12'b100110001101;
		if(({row_reg, col_reg}==14'b11000110101111)) color_data = 12'b101110101100;
		if(({row_reg, col_reg}==14'b11000110110000)) color_data = 12'b110010111011;
		if(({row_reg, col_reg}>=14'b11000110110001) && ({row_reg, col_reg}<14'b11000110110101)) color_data = 12'b101110101011;
		if(({row_reg, col_reg}==14'b11000110110101)) color_data = 12'b101010001001;
		if(({row_reg, col_reg}==14'b11000110110110)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}>=14'b11000110110111) && ({row_reg, col_reg}<14'b11000110111001)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}>=14'b11000110111001) && ({row_reg, col_reg}<14'b11000110111011)) color_data = 12'b011001000100;
		if(({row_reg, col_reg}==14'b11000110111011)) color_data = 12'b010101000100;
		if(({row_reg, col_reg}==14'b11000110111100)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==14'b11000110111101)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}==14'b11000110111110)) color_data = 12'b010100110011;
		if(({row_reg, col_reg}==14'b11000110111111)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}==14'b11000111000000)) color_data = 12'b010100110011;
		if(({row_reg, col_reg}==14'b11000111000001)) color_data = 12'b010000100011;
		if(({row_reg, col_reg}==14'b11000111000010)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}>=14'b11000111000011) && ({row_reg, col_reg}<14'b11000111000101)) color_data = 12'b001100010001;
		if(({row_reg, col_reg}>=14'b11000111000101) && ({row_reg, col_reg}<14'b11000111001100)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}>=14'b11000111001100) && ({row_reg, col_reg}<14'b11000111001110)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}>=14'b11000111001110) && ({row_reg, col_reg}<14'b11000111010000)) color_data = 12'b001100010001;
		if(({row_reg, col_reg}==14'b11000111010000)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==14'b11000111010001)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}==14'b11000111010010)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==14'b11000111010011)) color_data = 12'b001100010001;
		if(({row_reg, col_reg}==14'b11000111010100)) color_data = 12'b010000010001;
		if(({row_reg, col_reg}==14'b11000111010101)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}==14'b11000111010110)) color_data = 12'b010000100011;
		if(({row_reg, col_reg}>=14'b11000111010111) && ({row_reg, col_reg}<14'b11000111011101)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}==14'b11000111011101)) color_data = 12'b010000100011;
		if(({row_reg, col_reg}==14'b11000111011110)) color_data = 12'b010000100100;
		if(({row_reg, col_reg}==14'b11000111011111)) color_data = 12'b000100000100;
		if(({row_reg, col_reg}==14'b11000111100000)) color_data = 12'b000000001100;
		if(({row_reg, col_reg}==14'b11000111100001)) color_data = 12'b000000001101;
		if(({row_reg, col_reg}==14'b11000111100010)) color_data = 12'b000000001110;

		if(({row_reg, col_reg}>=14'b11000111100011) && ({row_reg, col_reg}<14'b11001000010000)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==14'b11001000010000)) color_data = 12'b000000001110;
		if(({row_reg, col_reg}==14'b11001000010001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==14'b11001000010010)) color_data = 12'b000000001110;
		if(({row_reg, col_reg}==14'b11001000010011)) color_data = 12'b000000001101;
		if(({row_reg, col_reg}==14'b11001000010100)) color_data = 12'b000000001011;
		if(({row_reg, col_reg}==14'b11001000010101)) color_data = 12'b000100001010;
		if(({row_reg, col_reg}==14'b11001000010110)) color_data = 12'b001000011001;
		if(({row_reg, col_reg}==14'b11001000010111)) color_data = 12'b001100011001;
		if(({row_reg, col_reg}==14'b11001000011000)) color_data = 12'b001100101000;
		if(({row_reg, col_reg}==14'b11001000011001)) color_data = 12'b010100111001;
		if(({row_reg, col_reg}==14'b11001000011010)) color_data = 12'b011001001001;
		if(({row_reg, col_reg}==14'b11001000011011)) color_data = 12'b001100101000;
		if(({row_reg, col_reg}==14'b11001000011100)) color_data = 12'b000100001000;
		if(({row_reg, col_reg}==14'b11001000011101)) color_data = 12'b000000001010;
		if(({row_reg, col_reg}==14'b11001000011110)) color_data = 12'b000000001100;
		if(({row_reg, col_reg}==14'b11001000011111)) color_data = 12'b000000001101;
		if(({row_reg, col_reg}==14'b11001000100000)) color_data = 12'b000000001110;
		if(({row_reg, col_reg}>=14'b11001000100001) && ({row_reg, col_reg}<14'b11001000101011)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==14'b11001000101011)) color_data = 12'b000000001101;
		if(({row_reg, col_reg}==14'b11001000101100)) color_data = 12'b001000101100;
		if(({row_reg, col_reg}==14'b11001000101101)) color_data = 12'b011001101100;
		if(({row_reg, col_reg}==14'b11001000101110)) color_data = 12'b101010011100;
		if(({row_reg, col_reg}>=14'b11001000101111) && ({row_reg, col_reg}<14'b11001000110011)) color_data = 12'b101110101011;
		if(({row_reg, col_reg}==14'b11001000110011)) color_data = 12'b110010101011;
		if(({row_reg, col_reg}==14'b11001000110100)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==14'b11001000110101)) color_data = 12'b100101111000;
		if(({row_reg, col_reg}>=14'b11001000110110) && ({row_reg, col_reg}<14'b11001000111000)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==14'b11001000111000)) color_data = 12'b101010001001;
		if(({row_reg, col_reg}==14'b11001000111001)) color_data = 12'b010000100011;
		if(({row_reg, col_reg}==14'b11001000111010)) color_data = 12'b001000000000;
		if(({row_reg, col_reg}==14'b11001000111011)) color_data = 12'b001100010001;
		if(({row_reg, col_reg}>=14'b11001000111100) && ({row_reg, col_reg}<14'b11001000111110)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}==14'b11001000111110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=14'b11001000111111) && ({row_reg, col_reg}<14'b11001001000011)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}==14'b11001001000011)) color_data = 12'b001100010001;
		if(({row_reg, col_reg}==14'b11001001000100)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==14'b11001001000101)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}==14'b11001001000110)) color_data = 12'b010000110011;
		if(({row_reg, col_reg}>=14'b11001001000111) && ({row_reg, col_reg}<14'b11001001001010)) color_data = 12'b010100110011;
		if(({row_reg, col_reg}>=14'b11001001001010) && ({row_reg, col_reg}<14'b11001001001100)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}>=14'b11001001001100) && ({row_reg, col_reg}<14'b11001001010000)) color_data = 12'b001100010001;
		if(({row_reg, col_reg}==14'b11001001010000)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}==14'b11001001010001)) color_data = 12'b010000110011;
		if(({row_reg, col_reg}==14'b11001001010010)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}>=14'b11001001010011) && ({row_reg, col_reg}<14'b11001001010101)) color_data = 12'b001100010001;
		if(({row_reg, col_reg}==14'b11001001010101)) color_data = 12'b010000100011;
		if(({row_reg, col_reg}==14'b11001001010110)) color_data = 12'b010100100011;
		if(({row_reg, col_reg}==14'b11001001010111)) color_data = 12'b010000100011;
		if(({row_reg, col_reg}>=14'b11001001011000) && ({row_reg, col_reg}<14'b11001001011010)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}==14'b11001001011010)) color_data = 12'b010000100011;
		if(({row_reg, col_reg}==14'b11001001011011)) color_data = 12'b010100100011;
		if(({row_reg, col_reg}==14'b11001001011100)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}==14'b11001001011101)) color_data = 12'b010000110011;
		if(({row_reg, col_reg}==14'b11001001011110)) color_data = 12'b010000100100;
		if(({row_reg, col_reg}==14'b11001001011111)) color_data = 12'b000100000100;
		if(({row_reg, col_reg}==14'b11001001100000)) color_data = 12'b000000001100;
		if(({row_reg, col_reg}==14'b11001001100001)) color_data = 12'b000000001101;
		if(({row_reg, col_reg}==14'b11001001100010)) color_data = 12'b000000001110;

		if(({row_reg, col_reg}>=14'b11001001100011) && ({row_reg, col_reg}<14'b11001010010000)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==14'b11001010010000)) color_data = 12'b000000001101;
		if(({row_reg, col_reg}==14'b11001010010001)) color_data = 12'b000100001101;
		if(({row_reg, col_reg}==14'b11001010010010)) color_data = 12'b000100001100;
		if(({row_reg, col_reg}==14'b11001010010011)) color_data = 12'b000100001010;
		if(({row_reg, col_reg}==14'b11001010010100)) color_data = 12'b001000011001;
		if(({row_reg, col_reg}==14'b11001010010101)) color_data = 12'b001100101001;
		if(({row_reg, col_reg}==14'b11001010010110)) color_data = 12'b010000111001;
		if(({row_reg, col_reg}>=14'b11001010010111) && ({row_reg, col_reg}<14'b11001010011010)) color_data = 12'b010100111001;
		if(({row_reg, col_reg}==14'b11001010011010)) color_data = 12'b010000101001;
		if(({row_reg, col_reg}==14'b11001010011011)) color_data = 12'b001000011000;
		if(({row_reg, col_reg}==14'b11001010011100)) color_data = 12'b000000001010;
		if(({row_reg, col_reg}==14'b11001010011101)) color_data = 12'b000000001100;
		if(({row_reg, col_reg}==14'b11001010011110)) color_data = 12'b000000001110;
		if(({row_reg, col_reg}==14'b11001010011111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==14'b11001010100000)) color_data = 12'b000000001110;
		if(({row_reg, col_reg}>=14'b11001010100001) && ({row_reg, col_reg}<14'b11001010101010)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==14'b11001010101010)) color_data = 12'b000000001110;
		if(({row_reg, col_reg}==14'b11001010101011)) color_data = 12'b000100011101;
		if(({row_reg, col_reg}==14'b11001010101100)) color_data = 12'b010001001100;
		if(({row_reg, col_reg}==14'b11001010101101)) color_data = 12'b100010001101;
		if(({row_reg, col_reg}==14'b11001010101110)) color_data = 12'b101110101100;
		if(({row_reg, col_reg}==14'b11001010101111)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}>=14'b11001010110000) && ({row_reg, col_reg}<14'b11001010110010)) color_data = 12'b101110101011;
		if(({row_reg, col_reg}==14'b11001010110010)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==14'b11001010110011)) color_data = 12'b101010011010;
		if(({row_reg, col_reg}==14'b11001010110100)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}>=14'b11001010110101) && ({row_reg, col_reg}<14'b11001010110111)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==14'b11001010110111)) color_data = 12'b011101010110;
		if(({row_reg, col_reg}==14'b11001010111000)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==14'b11001010111001)) color_data = 12'b010100110011;
		if(({row_reg, col_reg}==14'b11001010111010)) color_data = 12'b001100010001;
		if(({row_reg, col_reg}>=14'b11001010111011) && ({row_reg, col_reg}<14'b11001011000011)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}>=14'b11001011000011) && ({row_reg, col_reg}<14'b11001011000101)) color_data = 12'b001100010001;
		if(({row_reg, col_reg}>=14'b11001011000101) && ({row_reg, col_reg}<14'b11001011001011)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}==14'b11001011001011)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}>=14'b11001011001100) && ({row_reg, col_reg}<14'b11001011001110)) color_data = 12'b001100010001;
		if(({row_reg, col_reg}==14'b11001011001110)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}>=14'b11001011001111) && ({row_reg, col_reg}<14'b11001011010001)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}==14'b11001011010001)) color_data = 12'b010000110011;
		if(({row_reg, col_reg}==14'b11001011010010)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}>=14'b11001011010011) && ({row_reg, col_reg}<14'b11001011010101)) color_data = 12'b001100010001;
		if(({row_reg, col_reg}>=14'b11001011010101) && ({row_reg, col_reg}<14'b11001011011011)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}==14'b11001011011011)) color_data = 12'b010100100010;
		if(({row_reg, col_reg}==14'b11001011011100)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}==14'b11001011011101)) color_data = 12'b010000100011;
		if(({row_reg, col_reg}==14'b11001011011110)) color_data = 12'b001100100100;
		if(({row_reg, col_reg}==14'b11001011011111)) color_data = 12'b000100000011;
		if(({row_reg, col_reg}==14'b11001011100000)) color_data = 12'b000000001011;
		if(({row_reg, col_reg}==14'b11001011100001)) color_data = 12'b000000001101;
		if(({row_reg, col_reg}==14'b11001011100010)) color_data = 12'b000000001110;

		if(({row_reg, col_reg}>=14'b11001011100011) && ({row_reg, col_reg}<14'b11001100001101)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=14'b11001100001101) && ({row_reg, col_reg}<14'b11001100010000)) color_data = 12'b000000001110;
		if(({row_reg, col_reg}==14'b11001100010000)) color_data = 12'b000000001010;
		if(({row_reg, col_reg}==14'b11001100010001)) color_data = 12'b000100001010;
		if(({row_reg, col_reg}==14'b11001100010010)) color_data = 12'b001000001010;
		if(({row_reg, col_reg}==14'b11001100010011)) color_data = 12'b001000011000;
		if(({row_reg, col_reg}==14'b11001100010100)) color_data = 12'b001100101000;
		if(({row_reg, col_reg}==14'b11001100010101)) color_data = 12'b010101001000;
		if(({row_reg, col_reg}==14'b11001100010110)) color_data = 12'b010100111000;
		if(({row_reg, col_reg}==14'b11001100010111)) color_data = 12'b001100101000;
		if(({row_reg, col_reg}==14'b11001100011000)) color_data = 12'b001100101001;
		if(({row_reg, col_reg}==14'b11001100011001)) color_data = 12'b001000011001;
		if(({row_reg, col_reg}==14'b11001100011010)) color_data = 12'b000100001001;
		if(({row_reg, col_reg}==14'b11001100011011)) color_data = 12'b000000001011;
		if(({row_reg, col_reg}==14'b11001100011100)) color_data = 12'b000100001101;
		if(({row_reg, col_reg}==14'b11001100011101)) color_data = 12'b000000001110;
		if(({row_reg, col_reg}>=14'b11001100011110) && ({row_reg, col_reg}<14'b11001100101010)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==14'b11001100101010)) color_data = 12'b000000001110;
		if(({row_reg, col_reg}==14'b11001100101011)) color_data = 12'b001100101101;
		if(({row_reg, col_reg}==14'b11001100101100)) color_data = 12'b011001101101;
		if(({row_reg, col_reg}==14'b11001100101101)) color_data = 12'b101010011101;
		if(({row_reg, col_reg}==14'b11001100101110)) color_data = 12'b101110101011;
		if(({row_reg, col_reg}==14'b11001100101111)) color_data = 12'b110010101010;
		if(({row_reg, col_reg}==14'b11001100110000)) color_data = 12'b110010111011;
		if(({row_reg, col_reg}==14'b11001100110001)) color_data = 12'b101110101011;
		if(({row_reg, col_reg}==14'b11001100110010)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}>=14'b11001100110011) && ({row_reg, col_reg}<14'b11001100110110)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==14'b11001100110110)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==14'b11001100110111)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==14'b11001100111000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=14'b11001100111001) && ({row_reg, col_reg}<14'b11001100111011)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}==14'b11001100111011)) color_data = 12'b010000110011;
		if(({row_reg, col_reg}>=14'b11001100111100) && ({row_reg, col_reg}<14'b11001100111110)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}==14'b11001100111110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==14'b11001100111111)) color_data = 12'b010100110011;
		if(({row_reg, col_reg}==14'b11001101000000)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}==14'b11001101000001)) color_data = 12'b010000110011;
		if(({row_reg, col_reg}==14'b11001101000010)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}>=14'b11001101000011) && ({row_reg, col_reg}<14'b11001101001110)) color_data = 12'b001100010001;
		if(({row_reg, col_reg}>=14'b11001101001110) && ({row_reg, col_reg}<14'b11001101010001)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}==14'b11001101010001)) color_data = 12'b010000110011;
		if(({row_reg, col_reg}==14'b11001101010010)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}>=14'b11001101010011) && ({row_reg, col_reg}<14'b11001101010111)) color_data = 12'b001100010001;
		if(({row_reg, col_reg}==14'b11001101010111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==14'b11001101011000)) color_data = 12'b001100010001;
		if(({row_reg, col_reg}>=14'b11001101011001) && ({row_reg, col_reg}<14'b11001101011011)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}==14'b11001101011011)) color_data = 12'b010000100011;
		if(({row_reg, col_reg}>=14'b11001101011100) && ({row_reg, col_reg}<14'b11001101011110)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}==14'b11001101011110)) color_data = 12'b001100100011;
		if(({row_reg, col_reg}==14'b11001101011111)) color_data = 12'b000100000011;
		if(({row_reg, col_reg}==14'b11001101100000)) color_data = 12'b000000001011;
		if(({row_reg, col_reg}==14'b11001101100001)) color_data = 12'b000000001101;
		if(({row_reg, col_reg}==14'b11001101100010)) color_data = 12'b000000001110;

		if(({row_reg, col_reg}>=14'b11001101100011) && ({row_reg, col_reg}<14'b11001110001011)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==14'b11001110001011)) color_data = 12'b000000001110;
		if(({row_reg, col_reg}==14'b11001110001100)) color_data = 12'b000000001101;
		if(({row_reg, col_reg}==14'b11001110001101)) color_data = 12'b000000001100;
		if(({row_reg, col_reg}==14'b11001110001110)) color_data = 12'b000100001100;
		if(({row_reg, col_reg}==14'b11001110001111)) color_data = 12'b000100001011;
		if(({row_reg, col_reg}==14'b11001110010000)) color_data = 12'b001000001000;
		if(({row_reg, col_reg}==14'b11001110010001)) color_data = 12'b010000101010;
		if(({row_reg, col_reg}==14'b11001110010010)) color_data = 12'b010101001011;
		if(({row_reg, col_reg}==14'b11001110010011)) color_data = 12'b010100111010;
		if(({row_reg, col_reg}==14'b11001110010100)) color_data = 12'b010100111000;
		if(({row_reg, col_reg}==14'b11001110010101)) color_data = 12'b010101001000;
		if(({row_reg, col_reg}==14'b11001110010110)) color_data = 12'b001100101000;
		if(({row_reg, col_reg}==14'b11001110010111)) color_data = 12'b000100000111;
		if(({row_reg, col_reg}==14'b11001110011000)) color_data = 12'b000100001001;
		if(({row_reg, col_reg}==14'b11001110011001)) color_data = 12'b000000001010;
		if(({row_reg, col_reg}==14'b11001110011010)) color_data = 12'b000000001011;
		if(({row_reg, col_reg}==14'b11001110011011)) color_data = 12'b000000001101;
		if(({row_reg, col_reg}==14'b11001110011100)) color_data = 12'b000000001110;
		if(({row_reg, col_reg}>=14'b11001110011101) && ({row_reg, col_reg}<14'b11001110101010)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==14'b11001110101010)) color_data = 12'b000100001101;
		if(({row_reg, col_reg}==14'b11001110101011)) color_data = 12'b010001001100;
		if(({row_reg, col_reg}==14'b11001110101100)) color_data = 12'b100010001101;
		if(({row_reg, col_reg}==14'b11001110101101)) color_data = 12'b101110101100;
		if(({row_reg, col_reg}==14'b11001110101110)) color_data = 12'b101110101011;
		if(({row_reg, col_reg}==14'b11001110101111)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==14'b11001110110000)) color_data = 12'b101110101011;
		if(({row_reg, col_reg}==14'b11001110110001)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==14'b11001110110010)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==14'b11001110110011)) color_data = 12'b100101111000;
		if(({row_reg, col_reg}>=14'b11001110110100) && ({row_reg, col_reg}<14'b11001110110110)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==14'b11001110110110)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==14'b11001110110111)) color_data = 12'b001100010001;
		if(({row_reg, col_reg}==14'b11001110111000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=14'b11001110111001) && ({row_reg, col_reg}<14'b11001110111100)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}==14'b11001110111100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=14'b11001110111101) && ({row_reg, col_reg}<14'b11001111000010)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}==14'b11001111000010)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}>=14'b11001111000011) && ({row_reg, col_reg}<14'b11001111001010)) color_data = 12'b001100010001;
		if(({row_reg, col_reg}==14'b11001111001010)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=14'b11001111001011) && ({row_reg, col_reg}<14'b11001111001110)) color_data = 12'b001100010001;
		if(({row_reg, col_reg}>=14'b11001111001110) && ({row_reg, col_reg}<14'b11001111010001)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}==14'b11001111010001)) color_data = 12'b010000100011;
		if(({row_reg, col_reg}==14'b11001111010010)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}>=14'b11001111010011) && ({row_reg, col_reg}<14'b11001111011001)) color_data = 12'b001100010001;
		if(({row_reg, col_reg}==14'b11001111011001)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==14'b11001111011010)) color_data = 12'b010000100011;
		if(({row_reg, col_reg}==14'b11001111011011)) color_data = 12'b010100100011;
		if(({row_reg, col_reg}>=14'b11001111011100) && ({row_reg, col_reg}<14'b11001111011110)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}==14'b11001111011110)) color_data = 12'b001100100100;
		if(({row_reg, col_reg}==14'b11001111011111)) color_data = 12'b000100000011;
		if(({row_reg, col_reg}==14'b11001111100000)) color_data = 12'b000000001011;
		if(({row_reg, col_reg}==14'b11001111100001)) color_data = 12'b000000001101;
		if(({row_reg, col_reg}==14'b11001111100010)) color_data = 12'b000000001110;

		if(({row_reg, col_reg}>=14'b11001111100011) && ({row_reg, col_reg}<14'b11010000001010)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==14'b11010000001010)) color_data = 12'b000000001110;
		if(({row_reg, col_reg}==14'b11010000001011)) color_data = 12'b000000001100;
		if(({row_reg, col_reg}==14'b11010000001100)) color_data = 12'b000100001010;
		if(({row_reg, col_reg}==14'b11010000001101)) color_data = 12'b000100011001;
		if(({row_reg, col_reg}==14'b11010000001110)) color_data = 12'b001000011001;
		if(({row_reg, col_reg}==14'b11010000001111)) color_data = 12'b001100101001;
		if(({row_reg, col_reg}==14'b11010000010000)) color_data = 12'b010100111000;
		if(({row_reg, col_reg}==14'b11010000010001)) color_data = 12'b010100111001;
		if(({row_reg, col_reg}==14'b11010000010010)) color_data = 12'b010000111001;
		if(({row_reg, col_reg}>=14'b11010000010011) && ({row_reg, col_reg}<14'b11010000010101)) color_data = 12'b010000101000;
		if(({row_reg, col_reg}==14'b11010000010101)) color_data = 12'b001100011000;
		if(({row_reg, col_reg}==14'b11010000010110)) color_data = 12'b000100001001;
		if(({row_reg, col_reg}==14'b11010000010111)) color_data = 12'b000100001010;
		if(({row_reg, col_reg}==14'b11010000011000)) color_data = 12'b000000001100;
		if(({row_reg, col_reg}==14'b11010000011001)) color_data = 12'b000000001101;
		if(({row_reg, col_reg}==14'b11010000011010)) color_data = 12'b000000001110;
		if(({row_reg, col_reg}>=14'b11010000011011) && ({row_reg, col_reg}<14'b11010000101001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==14'b11010000101001)) color_data = 12'b000000001110;
		if(({row_reg, col_reg}==14'b11010000101010)) color_data = 12'b000100011100;
		if(({row_reg, col_reg}==14'b11010000101011)) color_data = 12'b011001101100;
		if(({row_reg, col_reg}==14'b11010000101100)) color_data = 12'b100110011100;
		if(({row_reg, col_reg}==14'b11010000101101)) color_data = 12'b101110101011;
		if(({row_reg, col_reg}==14'b11010000101110)) color_data = 12'b110010111011;
		if(({row_reg, col_reg}==14'b11010000101111)) color_data = 12'b110010101010;
		if(({row_reg, col_reg}==14'b11010000110000)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==14'b11010000110001)) color_data = 12'b110010101011;
		if(({row_reg, col_reg}==14'b11010000110010)) color_data = 12'b101010001001;
		if(({row_reg, col_reg}==14'b11010000110011)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==14'b11010000110100)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}>=14'b11010000110101) && ({row_reg, col_reg}<14'b11010000110111)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}>=14'b11010000110111) && ({row_reg, col_reg}<14'b11010000111001)) color_data = 12'b001100010001;
		if(({row_reg, col_reg}>=14'b11010000111001) && ({row_reg, col_reg}<14'b11010000111100)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}==14'b11010000111100)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=14'b11010000111101) && ({row_reg, col_reg}<14'b11010000111111)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}==14'b11010000111111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=14'b11010001000000) && ({row_reg, col_reg}<14'b11010001001100)) color_data = 12'b001100010001;
		if(({row_reg, col_reg}>=14'b11010001001100) && ({row_reg, col_reg}<14'b11010001010000)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}>=14'b11010001010000) && ({row_reg, col_reg}<14'b11010001011010)) color_data = 12'b001100010001;
		if(({row_reg, col_reg}>=14'b11010001011010) && ({row_reg, col_reg}<14'b11010001011110)) color_data = 12'b001100010010;
		if(({row_reg, col_reg}==14'b11010001011110)) color_data = 12'b001000010011;
		if(({row_reg, col_reg}==14'b11010001011111)) color_data = 12'b000100000011;
		if(({row_reg, col_reg}==14'b11010001100000)) color_data = 12'b000000001011;
		if(({row_reg, col_reg}==14'b11010001100001)) color_data = 12'b000000001101;
		if(({row_reg, col_reg}==14'b11010001100010)) color_data = 12'b000000001110;

		if(({row_reg, col_reg}>=14'b11010001100011) && ({row_reg, col_reg}<14'b11010010001001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==14'b11010010001001)) color_data = 12'b000000001110;
		if(({row_reg, col_reg}==14'b11010010001010)) color_data = 12'b000000001101;
		if(({row_reg, col_reg}==14'b11010010001011)) color_data = 12'b000100001011;
		if(({row_reg, col_reg}==14'b11010010001100)) color_data = 12'b001000101001;
		if(({row_reg, col_reg}==14'b11010010001101)) color_data = 12'b010000111001;
		if(({row_reg, col_reg}>=14'b11010010001110) && ({row_reg, col_reg}<14'b11010010010001)) color_data = 12'b010101001000;
		if(({row_reg, col_reg}==14'b11010010010001)) color_data = 12'b010000111000;
		if(({row_reg, col_reg}==14'b11010010010010)) color_data = 12'b001100011000;
		if(({row_reg, col_reg}==14'b11010010010011)) color_data = 12'b000100001000;
		if(({row_reg, col_reg}==14'b11010010010100)) color_data = 12'b000100001001;
		if(({row_reg, col_reg}==14'b11010010010101)) color_data = 12'b000000001010;
		if(({row_reg, col_reg}==14'b11010010010110)) color_data = 12'b000000001011;
		if(({row_reg, col_reg}==14'b11010010010111)) color_data = 12'b000000001101;
		if(({row_reg, col_reg}==14'b11010010011000)) color_data = 12'b000000001110;
		if(({row_reg, col_reg}>=14'b11010010011001) && ({row_reg, col_reg}<14'b11010010101001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==14'b11010010101001)) color_data = 12'b000000001101;
		if(({row_reg, col_reg}==14'b11010010101010)) color_data = 12'b010000111100;
		if(({row_reg, col_reg}==14'b11010010101011)) color_data = 12'b100001111100;
		if(({row_reg, col_reg}==14'b11010010101100)) color_data = 12'b101110101100;
		if(({row_reg, col_reg}==14'b11010010101101)) color_data = 12'b101110101011;
		if(({row_reg, col_reg}==14'b11010010101110)) color_data = 12'b110010101010;
		if(({row_reg, col_reg}==14'b11010010101111)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}>=14'b11010010110000) && ({row_reg, col_reg}<14'b11010010110010)) color_data = 12'b110010111011;
		if(({row_reg, col_reg}==14'b11010010110010)) color_data = 12'b101010001001;
		if(({row_reg, col_reg}==14'b11010010110011)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==14'b11010010110100)) color_data = 12'b011001010101;
		if(({row_reg, col_reg}==14'b11010010110101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=14'b11010010110110) && ({row_reg, col_reg}<14'b11010010111001)) color_data = 12'b001100010001;
		if(({row_reg, col_reg}==14'b11010010111001)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}==14'b11010010111010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==14'b11010010111011)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}>=14'b11010010111100) && ({row_reg, col_reg}<14'b11010010111110)) color_data = 12'b010100110010;
		if(({row_reg, col_reg}>=14'b11010010111110) && ({row_reg, col_reg}<14'b11010011000000)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}>=14'b11010011000000) && ({row_reg, col_reg}<14'b11010011001011)) color_data = 12'b001100010001;
		if(({row_reg, col_reg}==14'b11010011001011)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==14'b11010011001100)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}>=14'b11010011001101) && ({row_reg, col_reg}<14'b11010011010000)) color_data = 12'b010000110011;
		if(({row_reg, col_reg}>=14'b11010011010000) && ({row_reg, col_reg}<14'b11010011011010)) color_data = 12'b001100010001;
		if(({row_reg, col_reg}>=14'b11010011011010) && ({row_reg, col_reg}<14'b11010011011100)) color_data = 12'b001100010010;
		if(({row_reg, col_reg}>=14'b11010011011100) && ({row_reg, col_reg}<14'b11010011011110)) color_data = 12'b001100010001;
		if(({row_reg, col_reg}==14'b11010011011110)) color_data = 12'b001000010011;
		if(({row_reg, col_reg}==14'b11010011011111)) color_data = 12'b000000000011;
		if(({row_reg, col_reg}==14'b11010011100000)) color_data = 12'b000000001011;
		if(({row_reg, col_reg}==14'b11010011100001)) color_data = 12'b000000001101;
		if(({row_reg, col_reg}==14'b11010011100010)) color_data = 12'b000000001110;

		if(({row_reg, col_reg}>=14'b11010011100011) && ({row_reg, col_reg}<14'b11010100001001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==14'b11010100001001)) color_data = 12'b000000001110;
		if(({row_reg, col_reg}==14'b11010100001010)) color_data = 12'b000000001100;
		if(({row_reg, col_reg}==14'b11010100001011)) color_data = 12'b000100001010;
		if(({row_reg, col_reg}==14'b11010100001100)) color_data = 12'b001000011000;
		if(({row_reg, col_reg}==14'b11010100001101)) color_data = 12'b010000111000;
		if(({row_reg, col_reg}==14'b11010100001110)) color_data = 12'b010000110111;
		if(({row_reg, col_reg}==14'b11010100001111)) color_data = 12'b010000110110;
		if(({row_reg, col_reg}==14'b11010100010000)) color_data = 12'b010000111000;
		if(({row_reg, col_reg}==14'b11010100010001)) color_data = 12'b001100101001;
		if(({row_reg, col_reg}==14'b11010100010010)) color_data = 12'b000100001001;
		if(({row_reg, col_reg}==14'b11010100010011)) color_data = 12'b000000001010;
		if(({row_reg, col_reg}==14'b11010100010100)) color_data = 12'b000000001011;
		if(({row_reg, col_reg}==14'b11010100010101)) color_data = 12'b000000001101;
		if(({row_reg, col_reg}==14'b11010100010110)) color_data = 12'b000000001110;
		if(({row_reg, col_reg}>=14'b11010100010111) && ({row_reg, col_reg}<14'b11010100101000)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==14'b11010100101000)) color_data = 12'b000000001110;
		if(({row_reg, col_reg}==14'b11010100101001)) color_data = 12'b001000101101;
		if(({row_reg, col_reg}==14'b11010100101010)) color_data = 12'b011001011100;
		if(({row_reg, col_reg}==14'b11010100101011)) color_data = 12'b100110011100;
		if(({row_reg, col_reg}==14'b11010100101100)) color_data = 12'b101110101011;
		if(({row_reg, col_reg}==14'b11010100101101)) color_data = 12'b110010101011;
		if(({row_reg, col_reg}>=14'b11010100101110) && ({row_reg, col_reg}<14'b11010100110000)) color_data = 12'b110010101010;
		if(({row_reg, col_reg}>=14'b11010100110000) && ({row_reg, col_reg}<14'b11010100110010)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==14'b11010100110010)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==14'b11010100110011)) color_data = 12'b101010001001;
		if(({row_reg, col_reg}==14'b11010100110100)) color_data = 12'b011101010101;
		if(({row_reg, col_reg}==14'b11010100110101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==14'b11010100110110)) color_data = 12'b001100010001;
		if(({row_reg, col_reg}>=14'b11010100110111) && ({row_reg, col_reg}<14'b11010100111010)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}==14'b11010100111010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==14'b11010100111011)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}==14'b11010100111100)) color_data = 12'b001100010001;
		if(({row_reg, col_reg}>=14'b11010100111101) && ({row_reg, col_reg}<14'b11010100111111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==14'b11010100111111)) color_data = 12'b001100010001;
		if(({row_reg, col_reg}==14'b11010101000000)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}==14'b11010101000001)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}>=14'b11010101000010) && ({row_reg, col_reg}<14'b11010101000100)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}==14'b11010101000100)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}>=14'b11010101000101) && ({row_reg, col_reg}<14'b11010101001100)) color_data = 12'b001100010001;
		if(({row_reg, col_reg}>=14'b11010101001100) && ({row_reg, col_reg}<14'b11010101001110)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==14'b11010101001110)) color_data = 12'b001100010001;
		if(({row_reg, col_reg}==14'b11010101001111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=14'b11010101010000) && ({row_reg, col_reg}<14'b11010101011100)) color_data = 12'b001100010001;
		if(({row_reg, col_reg}==14'b11010101011100)) color_data = 12'b001100010000;
		if(({row_reg, col_reg}==14'b11010101011101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==14'b11010101011110)) color_data = 12'b001000010011;
		if(({row_reg, col_reg}==14'b11010101011111)) color_data = 12'b000000000011;
		if(({row_reg, col_reg}==14'b11010101100000)) color_data = 12'b000000001100;
		if(({row_reg, col_reg}==14'b11010101100001)) color_data = 12'b000000001101;
		if(({row_reg, col_reg}==14'b11010101100010)) color_data = 12'b000000001110;

		if(({row_reg, col_reg}>=14'b11010101100011) && ({row_reg, col_reg}<14'b11010110001001)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==14'b11010110001001)) color_data = 12'b000000001110;
		if(({row_reg, col_reg}==14'b11010110001010)) color_data = 12'b000000001101;
		if(({row_reg, col_reg}==14'b11010110001011)) color_data = 12'b000000001010;
		if(({row_reg, col_reg}==14'b11010110001100)) color_data = 12'b000000001000;
		if(({row_reg, col_reg}==14'b11010110001101)) color_data = 12'b000100000111;
		if(({row_reg, col_reg}>=14'b11010110001110) && ({row_reg, col_reg}<14'b11010110010000)) color_data = 12'b000100000110;
		if(({row_reg, col_reg}==14'b11010110010000)) color_data = 12'b000100001001;
		if(({row_reg, col_reg}==14'b11010110010001)) color_data = 12'b000000001001;
		if(({row_reg, col_reg}==14'b11010110010010)) color_data = 12'b000000001011;
		if(({row_reg, col_reg}==14'b11010110010011)) color_data = 12'b000000001101;
		if(({row_reg, col_reg}==14'b11010110010100)) color_data = 12'b000000001110;
		if(({row_reg, col_reg}>=14'b11010110010101) && ({row_reg, col_reg}<14'b11010110101000)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==14'b11010110101000)) color_data = 12'b000000001101;
		if(({row_reg, col_reg}==14'b11010110101001)) color_data = 12'b010001001101;
		if(({row_reg, col_reg}==14'b11010110101010)) color_data = 12'b100001111101;
		if(({row_reg, col_reg}==14'b11010110101011)) color_data = 12'b101010101100;
		if(({row_reg, col_reg}==14'b11010110101100)) color_data = 12'b101110101011;
		if(({row_reg, col_reg}>=14'b11010110101101) && ({row_reg, col_reg}<14'b11010110101111)) color_data = 12'b110010101011;
		if(({row_reg, col_reg}==14'b11010110101111)) color_data = 12'b110010111011;
		if(({row_reg, col_reg}==14'b11010110110000)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}>=14'b11010110110001) && ({row_reg, col_reg}<14'b11010110110011)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==14'b11010110110011)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==14'b11010110110100)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}>=14'b11010110110101) && ({row_reg, col_reg}<14'b11010110110111)) color_data = 12'b001100010001;
		if(({row_reg, col_reg}==14'b11010110110111)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}==14'b11010110111000)) color_data = 12'b010000110011;
		if(({row_reg, col_reg}==14'b11010110111001)) color_data = 12'b010100110011;
		if(({row_reg, col_reg}==14'b11010110111010)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==14'b11010110111011)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}==14'b11010110111100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=14'b11010110111101) && ({row_reg, col_reg}<14'b11010111000000)) color_data = 12'b001100010001;
		if(({row_reg, col_reg}>=14'b11010111000000) && ({row_reg, col_reg}<14'b11010111000010)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}>=14'b11010111000010) && ({row_reg, col_reg}<14'b11010111000100)) color_data = 12'b010100110011;
		if(({row_reg, col_reg}==14'b11010111000100)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}>=14'b11010111000101) && ({row_reg, col_reg}<14'b11010111001110)) color_data = 12'b001100010001;
		if(({row_reg, col_reg}==14'b11010111001110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=14'b11010111001111) && ({row_reg, col_reg}<14'b11010111010010)) color_data = 12'b001100010001;
		if(({row_reg, col_reg}==14'b11010111010010)) color_data = 12'b001100010010;
		if(({row_reg, col_reg}>=14'b11010111010011) && ({row_reg, col_reg}<14'b11010111011100)) color_data = 12'b001100010001;
		if(({row_reg, col_reg}==14'b11010111011100)) color_data = 12'b001100010000;
		if(({row_reg, col_reg}==14'b11010111011101)) color_data = 12'b001000100001;
		if(({row_reg, col_reg}==14'b11010111011110)) color_data = 12'b001000010011;
		if(({row_reg, col_reg}==14'b11010111011111)) color_data = 12'b000000000011;
		if(({row_reg, col_reg}==14'b11010111100000)) color_data = 12'b000000001100;
		if(({row_reg, col_reg}==14'b11010111100001)) color_data = 12'b000000001101;

		if(({row_reg, col_reg}>=14'b11010111100010) && ({row_reg, col_reg}<14'b11011000001010)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==14'b11011000001010)) color_data = 12'b000000001110;
		if(({row_reg, col_reg}==14'b11011000001011)) color_data = 12'b000000001100;
		if(({row_reg, col_reg}==14'b11011000001100)) color_data = 12'b000000001011;
		if(({row_reg, col_reg}>=14'b11011000001101) && ({row_reg, col_reg}<14'b11011000001111)) color_data = 12'b000000001010;
		if(({row_reg, col_reg}==14'b11011000001111)) color_data = 12'b000100001010;
		if(({row_reg, col_reg}==14'b11011000010000)) color_data = 12'b000000001011;
		if(({row_reg, col_reg}==14'b11011000010001)) color_data = 12'b000000001100;
		if(({row_reg, col_reg}==14'b11011000010010)) color_data = 12'b000000001110;
		if(({row_reg, col_reg}>=14'b11011000010011) && ({row_reg, col_reg}<14'b11011000100111)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==14'b11011000100111)) color_data = 12'b000000001110;
		if(({row_reg, col_reg}==14'b11011000101000)) color_data = 12'b000100011100;
		if(({row_reg, col_reg}==14'b11011000101001)) color_data = 12'b011001011101;
		if(({row_reg, col_reg}==14'b11011000101010)) color_data = 12'b100110011101;
		if(({row_reg, col_reg}==14'b11011000101011)) color_data = 12'b101110101100;
		if(({row_reg, col_reg}==14'b11011000101100)) color_data = 12'b110010101011;
		if(({row_reg, col_reg}==14'b11011000101101)) color_data = 12'b101110101011;
		if(({row_reg, col_reg}>=14'b11011000101110) && ({row_reg, col_reg}<14'b11011000110000)) color_data = 12'b101010011010;
		if(({row_reg, col_reg}>=14'b11011000110000) && ({row_reg, col_reg}<14'b11011000110010)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==14'b11011000110010)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==14'b11011000110011)) color_data = 12'b011101010101;
		if(({row_reg, col_reg}==14'b11011000110100)) color_data = 12'b010100110100;
		if(({row_reg, col_reg}==14'b11011000110101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==14'b11011000110110)) color_data = 12'b001100010001;
		if(({row_reg, col_reg}>=14'b11011000110111) && ({row_reg, col_reg}<14'b11011000111100)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}==14'b11011000111100)) color_data = 12'b001100010001;
		if(({row_reg, col_reg}==14'b11011000111101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==14'b11011000111110)) color_data = 12'b001100010001;
		if(({row_reg, col_reg}==14'b11011000111111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=14'b11011001000000) && ({row_reg, col_reg}<14'b11011001000100)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}==14'b11011001000100)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==14'b11011001000101)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}==14'b11011001000110)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}>=14'b11011001000111) && ({row_reg, col_reg}<14'b11011001011010)) color_data = 12'b001100010001;
		if(({row_reg, col_reg}>=14'b11011001011010) && ({row_reg, col_reg}<14'b11011001011101)) color_data = 12'b001100010000;
		if(({row_reg, col_reg}==14'b11011001011101)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==14'b11011001011110)) color_data = 12'b001000010011;
		if(({row_reg, col_reg}==14'b11011001011111)) color_data = 12'b000000000100;
		if(({row_reg, col_reg}==14'b11011001100000)) color_data = 12'b000000001100;
		if(({row_reg, col_reg}==14'b11011001100001)) color_data = 12'b000000001101;

		if(({row_reg, col_reg}>=14'b11011001100010) && ({row_reg, col_reg}<14'b11011010001011)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==14'b11011010001011)) color_data = 12'b000000001110;
		if(({row_reg, col_reg}>=14'b11011010001100) && ({row_reg, col_reg}<14'b11011010001111)) color_data = 12'b000000001101;
		if(({row_reg, col_reg}>=14'b11011010001111) && ({row_reg, col_reg}<14'b11011010010010)) color_data = 12'b000000001110;
		if(({row_reg, col_reg}>=14'b11011010010010) && ({row_reg, col_reg}<14'b11011010100110)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==14'b11011010100110)) color_data = 12'b000000001110;
		if(({row_reg, col_reg}==14'b11011010100111)) color_data = 12'b000000001101;
		if(({row_reg, col_reg}==14'b11011010101000)) color_data = 12'b001000101011;
		if(({row_reg, col_reg}==14'b11011010101001)) color_data = 12'b011101101100;
		if(({row_reg, col_reg}==14'b11011010101010)) color_data = 12'b101110101100;
		if(({row_reg, col_reg}==14'b11011010101011)) color_data = 12'b110010101100;
		if(({row_reg, col_reg}==14'b11011010101100)) color_data = 12'b110010101011;
		if(({row_reg, col_reg}==14'b11011010101101)) color_data = 12'b101110011011;
		if(({row_reg, col_reg}==14'b11011010101110)) color_data = 12'b100110001001;
		if(({row_reg, col_reg}==14'b11011010101111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=14'b11011010110000) && ({row_reg, col_reg}<14'b11011010110010)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==14'b11011010110010)) color_data = 12'b010100110011;
		if(({row_reg, col_reg}>=14'b11011010110011) && ({row_reg, col_reg}<14'b11011010110101)) color_data = 12'b001100010001;
		if(({row_reg, col_reg}==14'b11011010110101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==14'b11011010110110)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}>=14'b11011010110111) && ({row_reg, col_reg}<14'b11011010111001)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}>=14'b11011010111001) && ({row_reg, col_reg}<14'b11011010111111)) color_data = 12'b001100010001;
		if(({row_reg, col_reg}==14'b11011010111111)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=14'b11011011000000) && ({row_reg, col_reg}<14'b11011011000100)) color_data = 12'b001100010001;
		if(({row_reg, col_reg}==14'b11011011000100)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==14'b11011011000101)) color_data = 12'b010000110011;
		if(({row_reg, col_reg}==14'b11011011000110)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}>=14'b11011011000111) && ({row_reg, col_reg}<14'b11011011011010)) color_data = 12'b001100010001;
		if(({row_reg, col_reg}==14'b11011011011010)) color_data = 12'b001100010000;
		if(({row_reg, col_reg}>=14'b11011011011011) && ({row_reg, col_reg}<14'b11011011011101)) color_data = 12'b001100010001;
		if(({row_reg, col_reg}==14'b11011011011101)) color_data = 12'b001000010010;
		if(({row_reg, col_reg}==14'b11011011011110)) color_data = 12'b000100010101;
		if(({row_reg, col_reg}==14'b11011011011111)) color_data = 12'b000000000110;
		if(({row_reg, col_reg}==14'b11011011100000)) color_data = 12'b000000001101;
		if(({row_reg, col_reg}==14'b11011011100001)) color_data = 12'b000000001110;

		if(({row_reg, col_reg}>=14'b11011011100010) && ({row_reg, col_reg}<14'b11011100001100)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=14'b11011100001100) && ({row_reg, col_reg}<14'b11011100001110)) color_data = 12'b000000001110;
		if(({row_reg, col_reg}>=14'b11011100001110) && ({row_reg, col_reg}<14'b11011100010000)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==14'b11011100010000)) color_data = 12'b000000001110;
		if(({row_reg, col_reg}>=14'b11011100010001) && ({row_reg, col_reg}<14'b11011100100110)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==14'b11011100100110)) color_data = 12'b000000001110;
		if(({row_reg, col_reg}==14'b11011100100111)) color_data = 12'b000100011101;
		if(({row_reg, col_reg}==14'b11011100101000)) color_data = 12'b010101001100;
		if(({row_reg, col_reg}==14'b11011100101001)) color_data = 12'b100110011100;
		if(({row_reg, col_reg}==14'b11011100101010)) color_data = 12'b110010101100;
		if(({row_reg, col_reg}>=14'b11011100101011) && ({row_reg, col_reg}<14'b11011100101101)) color_data = 12'b110010101011;
		if(({row_reg, col_reg}==14'b11011100101101)) color_data = 12'b101010011010;
		if(({row_reg, col_reg}==14'b11011100101110)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==14'b11011100101111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=14'b11011100110000) && ({row_reg, col_reg}<14'b11011100110010)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==14'b11011100110010)) color_data = 12'b010000110011;
		if(({row_reg, col_reg}==14'b11011100110011)) color_data = 12'b001000000000;
		if(({row_reg, col_reg}>=14'b11011100110100) && ({row_reg, col_reg}<14'b11011100110111)) color_data = 12'b001100010001;
		if(({row_reg, col_reg}>=14'b11011100110111) && ({row_reg, col_reg}<14'b11011100111001)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}>=14'b11011100111001) && ({row_reg, col_reg}<14'b11011101000101)) color_data = 12'b001100010001;
		if(({row_reg, col_reg}>=14'b11011101000101) && ({row_reg, col_reg}<14'b11011101000111)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}>=14'b11011101000111) && ({row_reg, col_reg}<14'b11011101011100)) color_data = 12'b001100010001;
		if(({row_reg, col_reg}==14'b11011101011100)) color_data = 12'b001000010010;
		if(({row_reg, col_reg}==14'b11011101011101)) color_data = 12'b001000000011;
		if(({row_reg, col_reg}==14'b11011101011110)) color_data = 12'b000100000110;
		if(({row_reg, col_reg}==14'b11011101011111)) color_data = 12'b000000001000;
		if(({row_reg, col_reg}==14'b11011101100000)) color_data = 12'b000000001101;
		if(({row_reg, col_reg}==14'b11011101100001)) color_data = 12'b000000001110;

		if(({row_reg, col_reg}>=14'b11011101100010) && ({row_reg, col_reg}<14'b11011110010000)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==14'b11011110010000)) color_data = 12'b000000001110;
		if(({row_reg, col_reg}>=14'b11011110010001) && ({row_reg, col_reg}<14'b11011110100110)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==14'b11011110100110)) color_data = 12'b000100011110;
		if(({row_reg, col_reg}==14'b11011110100111)) color_data = 12'b001100111101;
		if(({row_reg, col_reg}==14'b11011110101000)) color_data = 12'b011101111101;
		if(({row_reg, col_reg}==14'b11011110101001)) color_data = 12'b101110101101;
		if(({row_reg, col_reg}==14'b11011110101010)) color_data = 12'b110010101011;
		if(({row_reg, col_reg}>=14'b11011110101011) && ({row_reg, col_reg}<14'b11011110101101)) color_data = 12'b101010001001;
		if(({row_reg, col_reg}==14'b11011110101101)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==14'b11011110101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==14'b11011110101111)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==14'b11011110110000)) color_data = 12'b100101110111;
		if(({row_reg, col_reg}==14'b11011110110001)) color_data = 12'b101010001000;
		if(({row_reg, col_reg}==14'b11011110110010)) color_data = 12'b010101000100;
		if(({row_reg, col_reg}==14'b11011110110011)) color_data = 12'b001000000000;
		if(({row_reg, col_reg}==14'b11011110110100)) color_data = 12'b001100010010;
		if(({row_reg, col_reg}>=14'b11011110110101) && ({row_reg, col_reg}<14'b11011110111101)) color_data = 12'b001100010001;
		if(({row_reg, col_reg}>=14'b11011110111101) && ({row_reg, col_reg}<14'b11011111000000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=14'b11011111000000) && ({row_reg, col_reg}<14'b11011111001110)) color_data = 12'b001100010001;
		if(({row_reg, col_reg}==14'b11011111001110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==14'b11011111001111)) color_data = 12'b001100010001;
		if(({row_reg, col_reg}==14'b11011111010000)) color_data = 12'b001100010000;
		if(({row_reg, col_reg}>=14'b11011111010001) && ({row_reg, col_reg}<14'b11011111011100)) color_data = 12'b001100010001;
		if(({row_reg, col_reg}==14'b11011111011100)) color_data = 12'b001000010010;
		if(({row_reg, col_reg}==14'b11011111011101)) color_data = 12'b000100000100;
		if(({row_reg, col_reg}==14'b11011111011110)) color_data = 12'b000100000111;
		if(({row_reg, col_reg}==14'b11011111011111)) color_data = 12'b000100001010;
		if(({row_reg, col_reg}==14'b11011111100000)) color_data = 12'b000000001101;
		if(({row_reg, col_reg}==14'b11011111100001)) color_data = 12'b000000001110;

		if(({row_reg, col_reg}>=14'b11011111100010) && ({row_reg, col_reg}<14'b11100000100101)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==14'b11100000100101)) color_data = 12'b000000001110;
		if(({row_reg, col_reg}==14'b11100000100110)) color_data = 12'b001000011100;
		if(({row_reg, col_reg}==14'b11100000100111)) color_data = 12'b011001101100;
		if(({row_reg, col_reg}==14'b11100000101000)) color_data = 12'b101010011100;
		if(({row_reg, col_reg}==14'b11100000101001)) color_data = 12'b101110101100;
		if(({row_reg, col_reg}==14'b11100000101010)) color_data = 12'b110010111100;
		if(({row_reg, col_reg}==14'b11100000101011)) color_data = 12'b101010011010;
		if(({row_reg, col_reg}==14'b11100000101100)) color_data = 12'b100110001001;
		if(({row_reg, col_reg}==14'b11100000101101)) color_data = 12'b100101111000;
		if(({row_reg, col_reg}==14'b11100000101110)) color_data = 12'b101010001001;
		if(({row_reg, col_reg}==14'b11100000101111)) color_data = 12'b100101111000;
		if(({row_reg, col_reg}>=14'b11100000110000) && ({row_reg, col_reg}<14'b11100000110010)) color_data = 12'b101010001000;
		if(({row_reg, col_reg}==14'b11100000110010)) color_data = 12'b010100110100;
		if(({row_reg, col_reg}==14'b11100000110011)) color_data = 12'b001000000001;
		if(({row_reg, col_reg}>=14'b11100000110100) && ({row_reg, col_reg}<14'b11100000110110)) color_data = 12'b001100010010;
		if(({row_reg, col_reg}==14'b11100000110110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==14'b11100000110111)) color_data = 12'b001100010010;
		if(({row_reg, col_reg}>=14'b11100000111000) && ({row_reg, col_reg}<14'b11100001001000)) color_data = 12'b001100010001;
		if(({row_reg, col_reg}==14'b11100001001000)) color_data = 12'b001100010010;
		if(({row_reg, col_reg}>=14'b11100001001001) && ({row_reg, col_reg}<14'b11100001010110)) color_data = 12'b001100010001;
		if(({row_reg, col_reg}==14'b11100001010110)) color_data = 12'b001100010000;
		if(({row_reg, col_reg}>=14'b11100001010111) && ({row_reg, col_reg}<14'b11100001011001)) color_data = 12'b001100010001;
		if(({row_reg, col_reg}==14'b11100001011001)) color_data = 12'b001100010010;
		if(({row_reg, col_reg}==14'b11100001011010)) color_data = 12'b001100010001;
		if(({row_reg, col_reg}==14'b11100001011011)) color_data = 12'b001100010010;
		if(({row_reg, col_reg}==14'b11100001011100)) color_data = 12'b001000010010;
		if(({row_reg, col_reg}==14'b11100001011101)) color_data = 12'b000100000101;
		if(({row_reg, col_reg}==14'b11100001011110)) color_data = 12'b000000001010;
		if(({row_reg, col_reg}==14'b11100001011111)) color_data = 12'b000000001110;

		if(({row_reg, col_reg}>=14'b11100001100000) && ({row_reg, col_reg}<14'b11100010100101)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==14'b11100010100101)) color_data = 12'b000000001101;
		if(({row_reg, col_reg}==14'b11100010100110)) color_data = 12'b001100111100;
		if(({row_reg, col_reg}==14'b11100010100111)) color_data = 12'b100001111101;
		if(({row_reg, col_reg}==14'b11100010101000)) color_data = 12'b101110101100;
		if(({row_reg, col_reg}==14'b11100010101001)) color_data = 12'b101010011010;
		if(({row_reg, col_reg}==14'b11100010101010)) color_data = 12'b100110001001;
		if(({row_reg, col_reg}>=14'b11100010101011) && ({row_reg, col_reg}<14'b11100010101101)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==14'b11100010101101)) color_data = 12'b100101110111;
		if(({row_reg, col_reg}==14'b11100010101110)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==14'b11100010101111)) color_data = 12'b100101110111;
		if(({row_reg, col_reg}==14'b11100010110000)) color_data = 12'b010101000100;
		if(({row_reg, col_reg}==14'b11100010110001)) color_data = 12'b010100110011;
		if(({row_reg, col_reg}==14'b11100010110010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=14'b11100010110011) && ({row_reg, col_reg}<14'b11100011010010)) color_data = 12'b001100010001;
		if(({row_reg, col_reg}==14'b11100011010010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=14'b11100011010011) && ({row_reg, col_reg}<14'b11100011010101)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}>=14'b11100011010101) && ({row_reg, col_reg}<14'b11100011010111)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}>=14'b11100011010111) && ({row_reg, col_reg}<14'b11100011011001)) color_data = 12'b001100010001;
		if(({row_reg, col_reg}>=14'b11100011011001) && ({row_reg, col_reg}<14'b11100011011100)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}==14'b11100011011100)) color_data = 12'b001000010010;
		if(({row_reg, col_reg}==14'b11100011011101)) color_data = 12'b000000000100;
		if(({row_reg, col_reg}==14'b11100011011110)) color_data = 12'b000000001010;
		if(({row_reg, col_reg}==14'b11100011011111)) color_data = 12'b000000001110;

		if(({row_reg, col_reg}>=14'b11100011100000) && ({row_reg, col_reg}<14'b11100100100100)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==14'b11100100100100)) color_data = 12'b000000001101;
		if(({row_reg, col_reg}==14'b11100100100101)) color_data = 12'b000100011100;
		if(({row_reg, col_reg}==14'b11100100100110)) color_data = 12'b010101011100;
		if(({row_reg, col_reg}==14'b11100100100111)) color_data = 12'b101010011101;
		if(({row_reg, col_reg}==14'b11100100101000)) color_data = 12'b101110111100;
		if(({row_reg, col_reg}>=14'b11100100101001) && ({row_reg, col_reg}<14'b11100100110000)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==14'b11100100110000)) color_data = 12'b001100010001;
		if(({row_reg, col_reg}==14'b11100100110001)) color_data = 12'b001000000000;
		if(({row_reg, col_reg}==14'b11100100110010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==14'b11100100110011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}>=14'b11100100110100) && ({row_reg, col_reg}<14'b11100100110111)) color_data = 12'b001100010001;
		if(({row_reg, col_reg}==14'b11100100110111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=14'b11100100111000) && ({row_reg, col_reg}<14'b11100101010000)) color_data = 12'b001100010001;
		if(({row_reg, col_reg}>=14'b11100101010000) && ({row_reg, col_reg}<14'b11100101010010)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==14'b11100101010010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==14'b11100101010011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}>=14'b11100101010100) && ({row_reg, col_reg}<14'b11100101010110)) color_data = 12'b010100110011;
		if(({row_reg, col_reg}==14'b11100101010110)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==14'b11100101010111)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==14'b11100101011000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==14'b11100101011001)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}==14'b11100101011010)) color_data = 12'b010100110011;
		if(({row_reg, col_reg}==14'b11100101011011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==14'b11100101011100)) color_data = 12'b001000010010;
		if(({row_reg, col_reg}==14'b11100101011101)) color_data = 12'b000000000100;
		if(({row_reg, col_reg}==14'b11100101011110)) color_data = 12'b000000001010;
		if(({row_reg, col_reg}==14'b11100101011111)) color_data = 12'b000000001110;

		if(({row_reg, col_reg}>=14'b11100101100000) && ({row_reg, col_reg}<14'b11100110100011)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==14'b11100110100011)) color_data = 12'b000000001110;
		if(({row_reg, col_reg}==14'b11100110100100)) color_data = 12'b000100011101;
		if(({row_reg, col_reg}==14'b11100110100101)) color_data = 12'b010001001101;
		if(({row_reg, col_reg}==14'b11100110100110)) color_data = 12'b100001111101;
		if(({row_reg, col_reg}==14'b11100110100111)) color_data = 12'b101110101100;
		if(({row_reg, col_reg}==14'b11100110101000)) color_data = 12'b101010011010;
		if(({row_reg, col_reg}==14'b11100110101001)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==14'b11100110101010)) color_data = 12'b101010001001;
		if(({row_reg, col_reg}==14'b11100110101011)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==14'b11100110101100)) color_data = 12'b011001010101;
		if(({row_reg, col_reg}==14'b11100110101101)) color_data = 12'b011001100101;
		if(({row_reg, col_reg}>=14'b11100110101110) && ({row_reg, col_reg}<14'b11100110110000)) color_data = 12'b011001010101;
		if(({row_reg, col_reg}==14'b11100110110000)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==14'b11100110110001)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}>=14'b11100110110010) && ({row_reg, col_reg}<14'b11100111010000)) color_data = 12'b001100010001;
		if(({row_reg, col_reg}>=14'b11100111010000) && ({row_reg, col_reg}<14'b11100111010011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==14'b11100111010011)) color_data = 12'b010000110011;
		if(({row_reg, col_reg}>=14'b11100111010100) && ({row_reg, col_reg}<14'b11100111010110)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==14'b11100111010110)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}>=14'b11100111010111) && ({row_reg, col_reg}<14'b11100111011001)) color_data = 12'b001100010001;
		if(({row_reg, col_reg}>=14'b11100111011001) && ({row_reg, col_reg}<14'b11100111011011)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==14'b11100111011011)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==14'b11100111011100)) color_data = 12'b001000010010;
		if(({row_reg, col_reg}==14'b11100111011101)) color_data = 12'b000000000101;
		if(({row_reg, col_reg}==14'b11100111011110)) color_data = 12'b000000001010;
		if(({row_reg, col_reg}==14'b11100111011111)) color_data = 12'b000000001110;

		if(({row_reg, col_reg}>=14'b11100111100000) && ({row_reg, col_reg}<14'b11101000100011)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==14'b11101000100011)) color_data = 12'b000000001101;
		if(({row_reg, col_reg}==14'b11101000100100)) color_data = 12'b001000011100;
		if(({row_reg, col_reg}==14'b11101000100101)) color_data = 12'b011001011101;
		if(({row_reg, col_reg}==14'b11101000100110)) color_data = 12'b100110001100;
		if(({row_reg, col_reg}==14'b11101000100111)) color_data = 12'b100110001001;
		if(({row_reg, col_reg}==14'b11101000101000)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==14'b11101000101001)) color_data = 12'b100101111000;
		if(({row_reg, col_reg}==14'b11101000101010)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==14'b11101000101011)) color_data = 12'b010100110100;
		if(({row_reg, col_reg}==14'b11101000101100)) color_data = 12'b000100000000;
		if(({row_reg, col_reg}==14'b11101000101101)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}>=14'b11101000101110) && ({row_reg, col_reg}<14'b11101000110000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}>=14'b11101000110000) && ({row_reg, col_reg}<14'b11101000110010)) color_data = 12'b010000110011;
		if(({row_reg, col_reg}==14'b11101000110010)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}>=14'b11101000110011) && ({row_reg, col_reg}<14'b11101000110101)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==14'b11101000110101)) color_data = 12'b001100010001;
		if(({row_reg, col_reg}>=14'b11101000110110) && ({row_reg, col_reg}<14'b11101000111000)) color_data = 12'b001100010010;
		if(({row_reg, col_reg}>=14'b11101000111000) && ({row_reg, col_reg}<14'b11101001001000)) color_data = 12'b001100010001;
		if(({row_reg, col_reg}==14'b11101001001000)) color_data = 12'b001100010010;
		if(({row_reg, col_reg}==14'b11101001001001)) color_data = 12'b001100010001;
		if(({row_reg, col_reg}>=14'b11101001001010) && ({row_reg, col_reg}<14'b11101001001100)) color_data = 12'b001100010010;
		if(({row_reg, col_reg}>=14'b11101001001100) && ({row_reg, col_reg}<14'b11101001010000)) color_data = 12'b001100010001;
		if(({row_reg, col_reg}==14'b11101001010000)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}==14'b11101001010001)) color_data = 12'b010100110011;
		if(({row_reg, col_reg}==14'b11101001010010)) color_data = 12'b010000110011;
		if(({row_reg, col_reg}==14'b11101001010011)) color_data = 12'b010100110100;
		if(({row_reg, col_reg}==14'b11101001010100)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==14'b11101001010101)) color_data = 12'b001100010010;
		if(({row_reg, col_reg}==14'b11101001010110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==14'b11101001010111)) color_data = 12'b001100010010;
		if(({row_reg, col_reg}==14'b11101001011000)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==14'b11101001011001)) color_data = 12'b001000000001;
		if(({row_reg, col_reg}>=14'b11101001011010) && ({row_reg, col_reg}<14'b11101001011100)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==14'b11101001011100)) color_data = 12'b000100000010;
		if(({row_reg, col_reg}==14'b11101001011101)) color_data = 12'b000000000110;
		if(({row_reg, col_reg}==14'b11101001011110)) color_data = 12'b000000001011;

		if(({row_reg, col_reg}>=14'b11101001011111) && ({row_reg, col_reg}<14'b11101010100011)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==14'b11101010100011)) color_data = 12'b000000001101;
		if(({row_reg, col_reg}==14'b11101010100100)) color_data = 12'b001100111101;
		if(({row_reg, col_reg}==14'b11101010100101)) color_data = 12'b100010001101;
		if(({row_reg, col_reg}==14'b11101010100110)) color_data = 12'b101010011011;
		if(({row_reg, col_reg}==14'b11101010100111)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==14'b11101010101000)) color_data = 12'b100001100110;
		if(({row_reg, col_reg}==14'b11101010101001)) color_data = 12'b101010001000;
		if(({row_reg, col_reg}==14'b11101010101010)) color_data = 12'b101010001001;
		if(({row_reg, col_reg}==14'b11101010101011)) color_data = 12'b011001010101;
		if(({row_reg, col_reg}==14'b11101010101100)) color_data = 12'b010000110011;
		if(({row_reg, col_reg}==14'b11101010101101)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}==14'b11101010101110)) color_data = 12'b001000000001;
		if(({row_reg, col_reg}==14'b11101010101111)) color_data = 12'b001000010010;
		if(({row_reg, col_reg}>=14'b11101010110000) && ({row_reg, col_reg}<14'b11101010110010)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}==14'b11101010110010)) color_data = 12'b001100010010;
		if(({row_reg, col_reg}==14'b11101010110011)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}==14'b11101010110100)) color_data = 12'b001100010010;
		if(({row_reg, col_reg}==14'b11101010110101)) color_data = 12'b001100010001;
		if(({row_reg, col_reg}==14'b11101010110110)) color_data = 12'b001100010010;
		if(({row_reg, col_reg}>=14'b11101010110111) && ({row_reg, col_reg}<14'b11101011001110)) color_data = 12'b001100010001;
		if(({row_reg, col_reg}>=14'b11101011001110) && ({row_reg, col_reg}<14'b11101011010000)) color_data = 12'b001100010010;
		if(({row_reg, col_reg}==14'b11101011010000)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}==14'b11101011010001)) color_data = 12'b010100110011;
		if(({row_reg, col_reg}>=14'b11101011010010) && ({row_reg, col_reg}<14'b11101011010100)) color_data = 12'b010000100011;
		if(({row_reg, col_reg}==14'b11101011010100)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==14'b11101011010101)) color_data = 12'b010000100011;
		if(({row_reg, col_reg}==14'b11101011010110)) color_data = 12'b001100010001;
		if(({row_reg, col_reg}==14'b11101011010111)) color_data = 12'b010000100011;
		if(({row_reg, col_reg}==14'b11101011011000)) color_data = 12'b010000110011;
		if(({row_reg, col_reg}==14'b11101011011001)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==14'b11101011011010)) color_data = 12'b010000110011;
		if(({row_reg, col_reg}==14'b11101011011011)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}==14'b11101011011100)) color_data = 12'b000100000010;
		if(({row_reg, col_reg}==14'b11101011011101)) color_data = 12'b000000000110;
		if(({row_reg, col_reg}==14'b11101011011110)) color_data = 12'b000000001011;

		if(({row_reg, col_reg}>=14'b11101011011111) && ({row_reg, col_reg}<14'b11101100100010)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==14'b11101100100010)) color_data = 12'b000000001110;
		if(({row_reg, col_reg}==14'b11101100100011)) color_data = 12'b000000001100;
		if(({row_reg, col_reg}==14'b11101100100100)) color_data = 12'b001100111011;
		if(({row_reg, col_reg}==14'b11101100100101)) color_data = 12'b011101111011;
		if(({row_reg, col_reg}==14'b11101100100110)) color_data = 12'b100001100111;
		if(({row_reg, col_reg}==14'b11101100100111)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==14'b11101100101000)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==14'b11101100101001)) color_data = 12'b101010001000;
		if(({row_reg, col_reg}==14'b11101100101010)) color_data = 12'b110010101011;
		if(({row_reg, col_reg}>=14'b11101100101011) && ({row_reg, col_reg}<14'b11101100101101)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==14'b11101100101101)) color_data = 12'b100101110111;
		if(({row_reg, col_reg}>=14'b11101100101110) && ({row_reg, col_reg}<14'b11101100110000)) color_data = 12'b001100010010;
		if(({row_reg, col_reg}>=14'b11101100110000) && ({row_reg, col_reg}<14'b11101100110010)) color_data = 12'b001100010001;
		if(({row_reg, col_reg}==14'b11101100110010)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==14'b11101100110011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==14'b11101100110100)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}>=14'b11101100110101) && ({row_reg, col_reg}<14'b11101101001110)) color_data = 12'b001100010001;
		if(({row_reg, col_reg}>=14'b11101101001110) && ({row_reg, col_reg}<14'b11101101010010)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}==14'b11101101010010)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==14'b11101101010011)) color_data = 12'b001100010001;
		if(({row_reg, col_reg}==14'b11101101010100)) color_data = 12'b010000110011;
		if(({row_reg, col_reg}>=14'b11101101010101) && ({row_reg, col_reg}<14'b11101101010111)) color_data = 12'b100101110111;
		if(({row_reg, col_reg}==14'b11101101010111)) color_data = 12'b101110101001;
		if(({row_reg, col_reg}==14'b11101101011000)) color_data = 12'b110010101010;
		if(({row_reg, col_reg}==14'b11101101011001)) color_data = 12'b101110101001;
		if(({row_reg, col_reg}==14'b11101101011010)) color_data = 12'b110010101010;
		if(({row_reg, col_reg}==14'b11101101011011)) color_data = 12'b100101110111;
		if(({row_reg, col_reg}==14'b11101101011100)) color_data = 12'b001100100100;
		if(({row_reg, col_reg}==14'b11101101011101)) color_data = 12'b000000000110;
		if(({row_reg, col_reg}==14'b11101101011110)) color_data = 12'b000000001011;
		if(({row_reg, col_reg}==14'b11101101011111)) color_data = 12'b000000001110;

		if(({row_reg, col_reg}>=14'b11101101100000) && ({row_reg, col_reg}<14'b11101110100010)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==14'b11101110100010)) color_data = 12'b000000001110;
		if(({row_reg, col_reg}==14'b11101110100011)) color_data = 12'b000100001100;
		if(({row_reg, col_reg}==14'b11101110100100)) color_data = 12'b010000111011;
		if(({row_reg, col_reg}==14'b11101110100101)) color_data = 12'b100001111011;
		if(({row_reg, col_reg}==14'b11101110100110)) color_data = 12'b011101100111;
		if(({row_reg, col_reg}>=14'b11101110100111) && ({row_reg, col_reg}<14'b11101110101001)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==14'b11101110101001)) color_data = 12'b101110011001;
		if(({row_reg, col_reg}==14'b11101110101010)) color_data = 12'b110010101011;
		if(({row_reg, col_reg}==14'b11101110101011)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==14'b11101110101100)) color_data = 12'b110110111100;
		if(({row_reg, col_reg}==14'b11101110101101)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==14'b11101110101110)) color_data = 12'b000100000001;
		if(({row_reg, col_reg}==14'b11101110101111)) color_data = 12'b001000010010;
		if(({row_reg, col_reg}==14'b11101110110000)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==14'b11101110110001)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==14'b11101110110010)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==14'b11101110110011)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==14'b11101110110100)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}>=14'b11101110110101) && ({row_reg, col_reg}<14'b11101110110111)) color_data = 12'b001100010000;
		if(({row_reg, col_reg}>=14'b11101110110111) && ({row_reg, col_reg}<14'b11101111001101)) color_data = 12'b001100010001;
		if(({row_reg, col_reg}==14'b11101111001101)) color_data = 12'b001100100001;
		if(({row_reg, col_reg}==14'b11101111001110)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}==14'b11101111001111)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==14'b11101111010000)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}==14'b11101111010001)) color_data = 12'b010000110010;
		if(({row_reg, col_reg}==14'b11101111010010)) color_data = 12'b010000100001;
		if(({row_reg, col_reg}==14'b11101111010011)) color_data = 12'b001000010000;
		if(({row_reg, col_reg}==14'b11101111010100)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==14'b11101111010101)) color_data = 12'b100110000111;
		if(({row_reg, col_reg}==14'b11101111010110)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==14'b11101111010111)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}>=14'b11101111011000) && ({row_reg, col_reg}<14'b11101111011010)) color_data = 12'b110010111010;
		if(({row_reg, col_reg}==14'b11101111011010)) color_data = 12'b110111001011;
		if(({row_reg, col_reg}==14'b11101111011011)) color_data = 12'b100101111000;
		if(({row_reg, col_reg}==14'b11101111011100)) color_data = 12'b000100000011;
		if(({row_reg, col_reg}==14'b11101111011101)) color_data = 12'b000000000110;
		if(({row_reg, col_reg}==14'b11101111011110)) color_data = 12'b000000001011;
		if(({row_reg, col_reg}==14'b11101111011111)) color_data = 12'b000000001110;

		if(({row_reg, col_reg}>=14'b11101111100000) && ({row_reg, col_reg}<14'b11110000100010)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==14'b11110000100010)) color_data = 12'b000000001110;
		if(({row_reg, col_reg}==14'b11110000100011)) color_data = 12'b000100001101;
		if(({row_reg, col_reg}==14'b11110000100100)) color_data = 12'b001000101010;
		if(({row_reg, col_reg}==14'b11110000100101)) color_data = 12'b001000100110;
		if(({row_reg, col_reg}==14'b11110000100110)) color_data = 12'b010000110101;
		if(({row_reg, col_reg}==14'b11110000100111)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==14'b11110000101000)) color_data = 12'b100001111000;
		if(({row_reg, col_reg}==14'b11110000101001)) color_data = 12'b100001111001;
		if(({row_reg, col_reg}>=14'b11110000101010) && ({row_reg, col_reg}<14'b11110000101101)) color_data = 12'b100110001010;
		if(({row_reg, col_reg}==14'b11110000101101)) color_data = 12'b100001111001;
		if(({row_reg, col_reg}==14'b11110000101110)) color_data = 12'b100001101000;
		if(({row_reg, col_reg}==14'b11110000101111)) color_data = 12'b011101101000;
		if(({row_reg, col_reg}>=14'b11110000110000) && ({row_reg, col_reg}<14'b11110000110010)) color_data = 12'b001100100011;
		if(({row_reg, col_reg}>=14'b11110000110010) && ({row_reg, col_reg}<14'b11110000111000)) color_data = 12'b001100010010;
		if(({row_reg, col_reg}>=14'b11110000111000) && ({row_reg, col_reg}<14'b11110001001011)) color_data = 12'b001000010010;
		if(({row_reg, col_reg}>=14'b11110001001011) && ({row_reg, col_reg}<14'b11110001001101)) color_data = 12'b001000010011;
		if(({row_reg, col_reg}==14'b11110001001101)) color_data = 12'b001100010011;
		if(({row_reg, col_reg}>=14'b11110001001110) && ({row_reg, col_reg}<14'b11110001010001)) color_data = 12'b001100100011;
		if(({row_reg, col_reg}==14'b11110001010001)) color_data = 12'b001100010010;
		if(({row_reg, col_reg}==14'b11110001010010)) color_data = 12'b001100100011;
		if(({row_reg, col_reg}==14'b11110001010011)) color_data = 12'b001000010010;
		if(({row_reg, col_reg}==14'b11110001010100)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}==14'b11110001010101)) color_data = 12'b100001111000;
		if(({row_reg, col_reg}>=14'b11110001010110) && ({row_reg, col_reg}<14'b11110001011010)) color_data = 12'b100110001010;
		if(({row_reg, col_reg}==14'b11110001011010)) color_data = 12'b100110001011;
		if(({row_reg, col_reg}==14'b11110001011011)) color_data = 12'b100001111010;
		if(({row_reg, col_reg}==14'b11110001011100)) color_data = 12'b010101001010;
		if(({row_reg, col_reg}==14'b11110001011101)) color_data = 12'b001000101010;
		if(({row_reg, col_reg}==14'b11110001011110)) color_data = 12'b000000001100;
		if(({row_reg, col_reg}==14'b11110001011111)) color_data = 12'b000000001110;

		if(({row_reg, col_reg}>=14'b11110001100000) && ({row_reg, col_reg}<14'b11110010100011)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==14'b11110010100011)) color_data = 12'b000000001101;
		if(({row_reg, col_reg}==14'b11110010100100)) color_data = 12'b000000001010;
		if(({row_reg, col_reg}==14'b11110010100101)) color_data = 12'b000000000110;
		if(({row_reg, col_reg}==14'b11110010100110)) color_data = 12'b001000010110;
		if(({row_reg, col_reg}==14'b11110010100111)) color_data = 12'b011001011001;
		if(({row_reg, col_reg}==14'b11110010101000)) color_data = 12'b011001011010;
		if(({row_reg, col_reg}==14'b11110010101001)) color_data = 12'b011001101010;
		if(({row_reg, col_reg}>=14'b11110010101010) && ({row_reg, col_reg}<14'b11110010101100)) color_data = 12'b011001101011;
		if(({row_reg, col_reg}==14'b11110010101100)) color_data = 12'b011001101010;
		if(({row_reg, col_reg}==14'b11110010101101)) color_data = 12'b011001011010;
		if(({row_reg, col_reg}==14'b11110010101110)) color_data = 12'b010101011010;
		if(({row_reg, col_reg}==14'b11110010101111)) color_data = 12'b010101001001;
		if(({row_reg, col_reg}==14'b11110010110000)) color_data = 12'b000000000101;
		if(({row_reg, col_reg}>=14'b11110010110001) && ({row_reg, col_reg}<14'b11110011010100)) color_data = 12'b000000000100;
		if(({row_reg, col_reg}==14'b11110011010100)) color_data = 12'b000100000110;
		if(({row_reg, col_reg}==14'b11110011010101)) color_data = 12'b010101001001;
		if(({row_reg, col_reg}>=14'b11110011010110) && ({row_reg, col_reg}<14'b11110011011010)) color_data = 12'b011001011011;
		if(({row_reg, col_reg}==14'b11110011011010)) color_data = 12'b011001011100;
		if(({row_reg, col_reg}==14'b11110011011011)) color_data = 12'b010101001100;
		if(({row_reg, col_reg}==14'b11110011011100)) color_data = 12'b001100111011;
		if(({row_reg, col_reg}==14'b11110011011101)) color_data = 12'b000100011100;
		if(({row_reg, col_reg}==14'b11110011011110)) color_data = 12'b000000001110;

		if(({row_reg, col_reg}>=14'b11110011011111) && ({row_reg, col_reg}<14'b11110100100100)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==14'b11110100100100)) color_data = 12'b000000001100;
		if(({row_reg, col_reg}==14'b11110100100101)) color_data = 12'b000000001010;
		if(({row_reg, col_reg}==14'b11110100100110)) color_data = 12'b000100001001;
		if(({row_reg, col_reg}==14'b11110100100111)) color_data = 12'b001000101010;
		if(({row_reg, col_reg}>=14'b11110100101000) && ({row_reg, col_reg}<14'b11110100101011)) color_data = 12'b001100101011;
		if(({row_reg, col_reg}>=14'b11110100101011) && ({row_reg, col_reg}<14'b11110100101111)) color_data = 12'b001000101011;
		if(({row_reg, col_reg}==14'b11110100101111)) color_data = 12'b001000011011;
		if(({row_reg, col_reg}>=14'b11110100110000) && ({row_reg, col_reg}<14'b11110101010101)) color_data = 12'b000000001001;
		if(({row_reg, col_reg}==14'b11110101010101)) color_data = 12'b001000011011;
		if(({row_reg, col_reg}>=14'b11110101010110) && ({row_reg, col_reg}<14'b11110101011100)) color_data = 12'b001000011100;
		if(({row_reg, col_reg}==14'b11110101011100)) color_data = 12'b000100011101;
		if(({row_reg, col_reg}==14'b11110101011101)) color_data = 12'b000000001110;

		if(({row_reg, col_reg}>=14'b11110101011110) && ({row_reg, col_reg}<14'b11110110100101)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}==14'b11110110100101)) color_data = 12'b000000001101;
		if(({row_reg, col_reg}>=14'b11110110100110) && ({row_reg, col_reg}<14'b11110110101001)) color_data = 12'b000000001100;
		if(({row_reg, col_reg}>=14'b11110110101001) && ({row_reg, col_reg}<14'b11110111010000)) color_data = 12'b000000001101;
		if(({row_reg, col_reg}==14'b11110111010000)) color_data = 12'b000000001110;
		if(({row_reg, col_reg}>=14'b11110111010001) && ({row_reg, col_reg}<14'b11110111010101)) color_data = 12'b000000001101;
		if(({row_reg, col_reg}==14'b11110111010101)) color_data = 12'b000000001110;
		if(({row_reg, col_reg}==14'b11110111010110)) color_data = 12'b000000001101;
		if(({row_reg, col_reg}>=14'b11110111010111) && ({row_reg, col_reg}<14'b11110111011001)) color_data = 12'b000000001110;
		if(({row_reg, col_reg}>=14'b11110111011001) && ({row_reg, col_reg}<14'b11110111011011)) color_data = 12'b000000001101;
		if(({row_reg, col_reg}>=14'b11110111011011) && ({row_reg, col_reg}<14'b11110111011101)) color_data = 12'b000000001110;

		if(({row_reg, col_reg}>=14'b11110111011101) && ({row_reg, col_reg}<14'b11111000100101)) color_data = 12'b000000001111;
		if(({row_reg, col_reg}>=14'b11111000100101) && ({row_reg, col_reg}<14'b11111000100111)) color_data = 12'b000000001110;




		if(({row_reg, col_reg}>=14'b11111000100111) && ({row_reg, col_reg}<=14'b11111111111111)) color_data = 12'b000000001111;
	end
endmodule